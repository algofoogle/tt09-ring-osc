magic
tech sky130A
magscale 1 2
timestamp 1731184872
<< viali >>
rect 6193 21641 6227 21675
rect 6745 21641 6779 21675
rect 7297 21641 7331 21675
rect 7849 21641 7883 21675
rect 8401 21641 8435 21675
rect 8953 21641 8987 21675
rect 9505 21641 9539 21675
rect 10057 21641 10091 21675
rect 10609 21641 10643 21675
rect 11161 21641 11195 21675
rect 11713 21641 11747 21675
rect 12265 21641 12299 21675
rect 12817 21641 12851 21675
rect 13553 21641 13587 21675
rect 13921 21641 13955 21675
rect 14473 21641 14507 21675
rect 15393 21641 15427 21675
rect 15669 21641 15703 21675
rect 16129 21641 16163 21675
rect 16773 21641 16807 21675
rect 16957 21641 16991 21675
rect 17601 21641 17635 21675
rect 18337 21641 18371 21675
rect 19901 21641 19935 21675
rect 24685 21641 24719 21675
rect 24869 21641 24903 21675
rect 26433 21641 26467 21675
rect 27077 21641 27111 21675
rect 19441 21573 19475 21607
rect 20545 21573 20579 21607
rect 22109 21573 22143 21607
rect 22201 21573 22235 21607
rect 23121 21573 23155 21607
rect 24961 21573 24995 21607
rect 26985 21573 27019 21607
rect 27353 21573 27387 21607
rect 29561 21573 29595 21607
rect 20177 21505 20211 21539
rect 25421 21505 25455 21539
rect 29101 21505 29135 21539
rect 15577 21437 15611 21471
rect 16589 21437 16623 21471
rect 17417 21437 17451 21471
rect 18521 21437 18555 21471
rect 19625 21437 19659 21471
rect 19717 21437 19751 21471
rect 20269 21437 20303 21471
rect 20361 21437 20395 21471
rect 20821 21437 20855 21471
rect 21005 21437 21039 21471
rect 21097 21437 21131 21471
rect 21281 21437 21315 21471
rect 21557 21437 21591 21471
rect 22385 21437 22419 21471
rect 22661 21437 22695 21471
rect 22753 21437 22787 21471
rect 23305 21437 23339 21471
rect 23673 21437 23707 21471
rect 24041 21437 24075 21471
rect 25145 21437 25179 21471
rect 25789 21437 25823 21471
rect 26249 21437 26283 21471
rect 26709 21437 26743 21471
rect 27261 21437 27295 21471
rect 27537 21437 27571 21471
rect 27813 21437 27847 21471
rect 27997 21437 28031 21471
rect 28089 21437 28123 21471
rect 28273 21437 28307 21471
rect 28365 21437 28399 21471
rect 28641 21437 28675 21471
rect 29009 21437 29043 21471
rect 29469 21437 29503 21471
rect 29745 21437 29779 21471
rect 20729 21369 20763 21403
rect 21833 21369 21867 21403
rect 23857 21369 23891 21403
rect 24501 21369 24535 21403
rect 25605 21369 25639 21403
rect 25973 21369 26007 21403
rect 26617 21369 26651 21403
rect 26801 21369 26835 21403
rect 21465 21301 21499 21335
rect 21741 21301 21775 21335
rect 21925 21301 21959 21335
rect 22477 21301 22511 21335
rect 22937 21301 22971 21335
rect 23397 21301 23431 21335
rect 23489 21301 23523 21335
rect 24133 21301 24167 21335
rect 24225 21301 24259 21335
rect 24409 21301 24443 21335
rect 24701 21301 24735 21335
rect 25697 21301 25731 21335
rect 26065 21301 26099 21335
rect 27721 21301 27755 21335
rect 28457 21301 28491 21335
rect 29377 21301 29411 21335
rect 15393 21097 15427 21131
rect 21373 21097 21407 21131
rect 21741 21097 21775 21131
rect 23673 21097 23707 21131
rect 23857 21097 23891 21131
rect 25145 21097 25179 21131
rect 26065 21097 26099 21131
rect 28457 21097 28491 21131
rect 29929 21097 29963 21131
rect 17601 21029 17635 21063
rect 27997 21029 28031 21063
rect 29377 21029 29411 21063
rect 12357 20961 12391 20995
rect 12449 20961 12483 20995
rect 12633 20961 12667 20995
rect 12725 20961 12759 20995
rect 12909 20961 12943 20995
rect 13001 20961 13035 20995
rect 13185 20961 13219 20995
rect 13277 20961 13311 20995
rect 13553 20961 13587 20995
rect 13645 20961 13679 20995
rect 13921 20961 13955 20995
rect 14013 20961 14047 20995
rect 14289 20961 14323 20995
rect 14933 20961 14967 20995
rect 15117 20961 15151 20995
rect 15209 20961 15243 20995
rect 15301 20961 15335 20995
rect 16589 20961 16623 20995
rect 16773 20961 16807 20995
rect 16865 20961 16899 20995
rect 17049 20961 17083 20995
rect 17141 20961 17175 20995
rect 17325 20961 17359 20995
rect 17417 20961 17451 20995
rect 17509 20961 17543 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 18889 20961 18923 20995
rect 19073 20961 19107 20995
rect 19165 20961 19199 20995
rect 19349 20961 19383 20995
rect 19441 20961 19475 20995
rect 19625 20961 19659 20995
rect 19717 20961 19751 20995
rect 19901 20961 19935 20995
rect 19993 20961 20027 20995
rect 20085 20961 20119 20995
rect 20177 20961 20211 20995
rect 20361 20961 20395 20995
rect 20453 20961 20487 20995
rect 20637 20961 20671 20995
rect 21465 20961 21499 20995
rect 21557 20961 21591 20995
rect 22017 20961 22051 20995
rect 22201 20961 22235 20995
rect 22293 20961 22327 20995
rect 22477 20961 22511 20995
rect 22569 20961 22603 20995
rect 22753 20961 22787 20995
rect 22845 20961 22879 20995
rect 23029 20961 23063 20995
rect 23121 20961 23155 20995
rect 23305 20961 23339 20995
rect 23397 20961 23431 20995
rect 23489 20961 23523 20995
rect 24041 20961 24075 20995
rect 24961 20961 24995 20995
rect 26249 20961 26283 20995
rect 26985 20961 27019 20995
rect 27169 20961 27203 20995
rect 27261 20961 27295 20995
rect 27445 20961 27479 20995
rect 27537 20961 27571 20995
rect 27721 20961 27755 20995
rect 27813 20961 27847 20995
rect 27905 20961 27939 20995
rect 28549 20961 28583 20995
rect 28825 20961 28859 20995
rect 29193 20961 29227 20995
rect 29285 20961 29319 20995
rect 29561 20961 29595 20995
rect 29653 20961 29687 20995
rect 29837 20961 29871 20995
rect 14381 20893 14415 20927
rect 21925 20893 21959 20927
rect 29101 20893 29135 20927
rect 28641 20825 28675 20859
rect 14841 20757 14875 20791
rect 16497 20757 16531 20791
rect 18521 20757 18555 20791
rect 20729 20757 20763 20791
rect 26893 20757 26927 20791
rect 12357 20553 12391 20587
rect 17509 20553 17543 20587
rect 19901 20553 19935 20587
rect 23305 20553 23339 20587
rect 29653 20553 29687 20587
rect 8493 20417 8527 20451
rect 12633 20417 12667 20451
rect 15117 20417 15151 20451
rect 17233 20417 17267 20451
rect 18429 20417 18463 20451
rect 19625 20417 19659 20451
rect 24501 20417 24535 20451
rect 1593 20349 1627 20383
rect 1869 20349 1903 20383
rect 3801 20349 3835 20383
rect 6469 20349 6503 20383
rect 6561 20349 6595 20383
rect 6745 20349 6779 20383
rect 6837 20349 6871 20383
rect 7021 20349 7055 20383
rect 7113 20349 7147 20383
rect 7297 20349 7331 20383
rect 7389 20349 7423 20383
rect 7573 20349 7607 20383
rect 8125 20349 8159 20383
rect 8401 20349 8435 20383
rect 11253 20349 11287 20383
rect 11345 20349 11379 20383
rect 11437 20349 11471 20383
rect 11621 20349 11655 20383
rect 12173 20349 12207 20383
rect 12265 20349 12299 20383
rect 12541 20349 12575 20383
rect 14657 20349 14691 20383
rect 14749 20349 14783 20383
rect 15025 20349 15059 20383
rect 16221 20349 16255 20383
rect 16405 20349 16439 20383
rect 16497 20349 16531 20383
rect 17325 20349 17359 20383
rect 17417 20349 17451 20383
rect 18521 20349 18555 20383
rect 18705 20349 18739 20383
rect 19717 20349 19751 20383
rect 19809 20349 19843 20383
rect 20821 20349 20855 20383
rect 20913 20349 20947 20383
rect 21097 20349 21131 20383
rect 21189 20349 21223 20383
rect 21373 20349 21407 20383
rect 23397 20349 23431 20383
rect 23581 20349 23615 20383
rect 23673 20349 23707 20383
rect 23949 20349 23983 20383
rect 24041 20349 24075 20383
rect 24225 20349 24259 20383
rect 24317 20349 24351 20383
rect 24409 20349 24443 20383
rect 26801 20349 26835 20383
rect 26985 20349 27019 20383
rect 27077 20349 27111 20383
rect 27261 20349 27295 20383
rect 27353 20349 27387 20383
rect 27445 20349 27479 20383
rect 29009 20349 29043 20383
rect 29101 20349 29135 20383
rect 29285 20349 29319 20383
rect 29377 20349 29411 20383
rect 29561 20349 29595 20383
rect 7665 20281 7699 20315
rect 11161 20281 11195 20315
rect 12081 20281 12115 20315
rect 14565 20281 14599 20315
rect 27537 20281 27571 20315
rect 1685 20213 1719 20247
rect 1961 20213 1995 20247
rect 3893 20213 3927 20247
rect 8033 20213 8067 20247
rect 11713 20213 11747 20247
rect 14841 20213 14875 20247
rect 16129 20213 16163 20247
rect 18797 20213 18831 20247
rect 21465 20213 21499 20247
rect 26709 20213 26743 20247
rect 1133 20009 1167 20043
rect 1409 20009 1443 20043
rect 3341 20009 3375 20043
rect 6469 20009 6503 20043
rect 11713 20009 11747 20043
rect 17693 20009 17727 20043
rect 19717 20009 19751 20043
rect 24225 20009 24259 20043
rect 2513 19941 2547 19975
rect 3617 19941 3651 19975
rect 4169 19941 4203 19975
rect 5273 19941 5307 19975
rect 6745 19941 6779 19975
rect 8861 19941 8895 19975
rect 11437 19941 11471 19975
rect 11989 19941 12023 19975
rect 13921 19941 13955 19975
rect 19165 19941 19199 19975
rect 20545 19941 20579 19975
rect 26157 19941 26191 19975
rect 28273 19941 28307 19975
rect 1225 19873 1259 19907
rect 1501 19873 1535 19907
rect 1777 19873 1811 19907
rect 1869 19873 1903 19907
rect 1961 19873 1995 19907
rect 2145 19873 2179 19907
rect 2605 19873 2639 19907
rect 2697 19873 2731 19907
rect 2789 19873 2823 19907
rect 2973 19873 3007 19907
rect 3065 19873 3099 19907
rect 3249 19873 3283 19907
rect 3709 19873 3743 19907
rect 3801 19873 3835 19907
rect 4261 19873 4295 19907
rect 4353 19873 4387 19907
rect 4445 19873 4479 19907
rect 4629 19873 4663 19907
rect 4721 19873 4755 19907
rect 4905 19873 4939 19907
rect 5365 19873 5399 19907
rect 5457 19873 5491 19907
rect 5549 19873 5583 19907
rect 6009 19873 6043 19907
rect 6561 19873 6595 19907
rect 6653 19873 6687 19907
rect 8125 19873 8159 19907
rect 8309 19873 8343 19907
rect 8401 19873 8435 19907
rect 8585 19873 8619 19907
rect 8677 19873 8711 19907
rect 8769 19873 8803 19907
rect 9597 19873 9631 19907
rect 10333 19873 10367 19907
rect 10609 19873 10643 19907
rect 11253 19873 11287 19907
rect 11345 19873 11379 19907
rect 11805 19873 11839 19907
rect 11897 19873 11931 19907
rect 12725 19873 12759 19907
rect 13185 19873 13219 19907
rect 13369 19873 13403 19907
rect 13461 19873 13495 19907
rect 13645 19873 13679 19907
rect 13737 19873 13771 19907
rect 14013 19873 14047 19907
rect 14197 19873 14231 19907
rect 14289 19873 14323 19907
rect 14381 19873 14415 19907
rect 15301 19873 15335 19907
rect 15485 19873 15519 19907
rect 15577 19873 15611 19907
rect 15761 19873 15795 19907
rect 15853 19873 15887 19907
rect 16129 19873 16163 19907
rect 17233 19873 17267 19907
rect 17325 19873 17359 19907
rect 17417 19873 17451 19907
rect 17601 19873 17635 19907
rect 18705 19873 18739 19907
rect 18889 19873 18923 19907
rect 18981 19873 19015 19907
rect 19073 19873 19107 19907
rect 19809 19873 19843 19907
rect 19993 19873 20027 19907
rect 20085 19873 20119 19907
rect 20177 19873 20211 19907
rect 20269 19873 20303 19907
rect 20453 19873 20487 19907
rect 21465 19873 21499 19907
rect 21557 19873 21591 19907
rect 21741 19873 21775 19907
rect 21833 19873 21867 19907
rect 22017 19873 22051 19907
rect 22109 19873 22143 19907
rect 22293 19873 22327 19907
rect 22385 19873 22419 19907
rect 22569 19873 22603 19907
rect 22661 19873 22695 19907
rect 22845 19873 22879 19907
rect 22937 19873 22971 19907
rect 23121 19873 23155 19907
rect 24317 19873 24351 19907
rect 24501 19873 24535 19907
rect 24593 19873 24627 19907
rect 24777 19873 24811 19907
rect 24869 19873 24903 19907
rect 25053 19873 25087 19907
rect 25145 19873 25179 19907
rect 25329 19873 25363 19907
rect 25421 19873 25455 19907
rect 25605 19873 25639 19907
rect 25697 19873 25731 19907
rect 25881 19873 25915 19907
rect 25973 19873 26007 19907
rect 26065 19873 26099 19907
rect 26617 19873 26651 19907
rect 26801 19873 26835 19907
rect 26893 19873 26927 19907
rect 27077 19873 27111 19907
rect 27169 19873 27203 19907
rect 27261 19873 27295 19907
rect 28365 19873 28399 19907
rect 28457 19873 28491 19907
rect 28549 19873 28583 19907
rect 28733 19873 28767 19907
rect 28825 19873 28859 19907
rect 29009 19873 29043 19907
rect 29101 19873 29135 19907
rect 29285 19873 29319 19907
rect 29377 19873 29411 19907
rect 29561 19873 29595 19907
rect 1685 19805 1719 19839
rect 6101 19805 6135 19839
rect 10701 19805 10735 19839
rect 14473 19805 14507 19839
rect 16221 19805 16255 19839
rect 17141 19805 17175 19839
rect 27353 19805 27387 19839
rect 11161 19737 11195 19771
rect 2237 19669 2271 19703
rect 3893 19669 3927 19703
rect 4997 19669 5031 19703
rect 8033 19669 8067 19703
rect 9689 19669 9723 19703
rect 10425 19669 10459 19703
rect 12633 19669 12667 19703
rect 13093 19669 13127 19703
rect 15209 19669 15243 19703
rect 18613 19669 18647 19703
rect 23213 19669 23247 19703
rect 26525 19669 26559 19703
rect 29653 19669 29687 19703
rect 2145 19465 2179 19499
rect 4445 19465 4479 19499
rect 8861 19465 8895 19499
rect 10149 19465 10183 19499
rect 10609 19465 10643 19499
rect 12817 19465 12851 19499
rect 17877 19465 17911 19499
rect 20177 19465 20211 19499
rect 25605 19465 25639 19499
rect 26617 19465 26651 19499
rect 28733 19465 28767 19499
rect 29101 19465 29135 19499
rect 23029 19397 23063 19431
rect 1501 19261 1535 19295
rect 1593 19261 1627 19295
rect 1777 19261 1811 19295
rect 1869 19261 1903 19295
rect 2053 19261 2087 19295
rect 2789 19261 2823 19295
rect 2881 19261 2915 19295
rect 3709 19261 3743 19295
rect 4353 19261 4387 19295
rect 5457 19261 5491 19295
rect 5549 19261 5583 19295
rect 7665 19261 7699 19295
rect 7849 19261 7883 19295
rect 7941 19261 7975 19295
rect 8125 19261 8159 19295
rect 8217 19261 8251 19295
rect 8401 19261 8435 19295
rect 8953 19261 8987 19295
rect 9137 19261 9171 19295
rect 9229 19261 9263 19295
rect 9321 19261 9355 19295
rect 9781 19261 9815 19295
rect 9873 19261 9907 19295
rect 10057 19261 10091 19295
rect 10517 19261 10551 19295
rect 12265 19261 12299 19295
rect 12357 19261 12391 19295
rect 12909 19261 12943 19295
rect 13001 19261 13035 19295
rect 13093 19261 13127 19295
rect 13553 19261 13587 19295
rect 15025 19261 15059 19295
rect 15209 19261 15243 19295
rect 15301 19261 15335 19295
rect 15669 19261 15703 19295
rect 15761 19261 15795 19295
rect 17141 19261 17175 19295
rect 17233 19261 17267 19295
rect 17325 19261 17359 19295
rect 17509 19261 17543 19295
rect 17601 19261 17635 19295
rect 17785 19261 17819 19295
rect 18889 19261 18923 19295
rect 19073 19261 19107 19295
rect 19165 19261 19199 19295
rect 19257 19261 19291 19295
rect 20269 19261 20303 19295
rect 20453 19261 20487 19295
rect 20545 19261 20579 19295
rect 20821 19261 20855 19295
rect 20913 19261 20947 19295
rect 22845 19261 22879 19295
rect 23121 19261 23155 19295
rect 23213 19261 23247 19295
rect 23489 19261 23523 19295
rect 25697 19261 25731 19295
rect 26709 19261 26743 19295
rect 28089 19261 28123 19295
rect 28181 19261 28215 19295
rect 28365 19261 28399 19295
rect 28457 19261 28491 19295
rect 28641 19261 28675 19295
rect 29193 19261 29227 19295
rect 8493 19193 8527 19227
rect 9413 19193 9447 19227
rect 12173 19193 12207 19227
rect 13645 19193 13679 19227
rect 15577 19193 15611 19227
rect 15853 19193 15887 19227
rect 17049 19193 17083 19227
rect 19349 19193 19383 19227
rect 20729 19193 20763 19227
rect 22753 19193 22787 19227
rect 23305 19193 23339 19227
rect 3801 19125 3835 19159
rect 7573 19125 7607 19159
rect 12449 19125 12483 19159
rect 14933 19125 14967 19159
rect 18797 19125 18831 19159
rect 21005 19125 21039 19159
rect 23581 19125 23615 19159
rect 1593 18921 1627 18955
rect 3525 18921 3559 18955
rect 9229 18921 9263 18955
rect 17785 18921 17819 18955
rect 20821 18921 20855 18955
rect 27997 18921 28031 18955
rect 2421 18853 2455 18887
rect 6193 18853 6227 18887
rect 8309 18853 8343 18887
rect 9873 18853 9907 18887
rect 13277 18853 13311 18887
rect 14565 18853 14599 18887
rect 19533 18853 19567 18887
rect 21373 18853 21407 18887
rect 23305 18853 23339 18887
rect 1685 18785 1719 18819
rect 1777 18785 1811 18819
rect 1869 18785 1903 18819
rect 2053 18785 2087 18819
rect 2145 18785 2179 18819
rect 2329 18785 2363 18819
rect 3433 18785 3467 18819
rect 3709 18785 3743 18819
rect 3801 18785 3835 18819
rect 3985 18785 4019 18819
rect 4077 18785 4111 18819
rect 4261 18785 4295 18819
rect 4353 18785 4387 18819
rect 4537 18785 4571 18819
rect 4629 18785 4663 18819
rect 4813 18785 4847 18819
rect 4905 18785 4939 18819
rect 5089 18785 5123 18819
rect 5181 18785 5215 18819
rect 5365 18785 5399 18819
rect 6009 18785 6043 18819
rect 6101 18785 6135 18819
rect 7297 18785 7331 18819
rect 7573 18785 7607 18819
rect 7757 18785 7791 18819
rect 7849 18785 7883 18819
rect 8033 18785 8067 18819
rect 8125 18785 8159 18819
rect 8217 18785 8251 18819
rect 9321 18785 9355 18819
rect 9505 18785 9539 18819
rect 9597 18785 9631 18819
rect 9965 18785 9999 18819
rect 10057 18785 10091 18819
rect 12265 18785 12299 18819
rect 12357 18785 12391 18819
rect 12817 18785 12851 18819
rect 13001 18785 13035 18819
rect 13093 18785 13127 18819
rect 13185 18785 13219 18819
rect 14657 18785 14691 18819
rect 14933 18785 14967 18819
rect 15117 18785 15151 18819
rect 15209 18785 15243 18819
rect 15393 18785 15427 18819
rect 15485 18785 15519 18819
rect 15577 18785 15611 18819
rect 16865 18785 16899 18819
rect 16957 18785 16991 18819
rect 17141 18785 17175 18819
rect 17233 18785 17267 18819
rect 17417 18785 17451 18819
rect 17509 18785 17543 18819
rect 17693 18785 17727 18819
rect 18797 18785 18831 18819
rect 19073 18785 19107 18819
rect 19257 18785 19291 18819
rect 19349 18785 19383 18819
rect 19441 18785 19475 18819
rect 20637 18785 20671 18819
rect 20913 18785 20947 18819
rect 21281 18785 21315 18819
rect 21557 18785 21591 18819
rect 21649 18785 21683 18819
rect 21833 18785 21867 18819
rect 23397 18785 23431 18819
rect 23489 18785 23523 18819
rect 23581 18785 23615 18819
rect 23765 18785 23799 18819
rect 23857 18785 23891 18819
rect 24041 18785 24075 18819
rect 24133 18785 24167 18819
rect 24317 18785 24351 18819
rect 24409 18785 24443 18819
rect 24593 18785 24627 18819
rect 24685 18785 24719 18819
rect 24869 18785 24903 18819
rect 24961 18785 24995 18819
rect 25145 18785 25179 18819
rect 25237 18785 25271 18819
rect 25421 18785 25455 18819
rect 25513 18785 25547 18819
rect 25697 18785 25731 18819
rect 28089 18785 28123 18819
rect 28273 18785 28307 18819
rect 28365 18785 28399 18819
rect 28457 18785 28491 18819
rect 28733 18785 28767 18819
rect 5457 18717 5491 18751
rect 7205 18717 7239 18751
rect 10149 18717 10183 18751
rect 12173 18717 12207 18751
rect 12449 18717 12483 18751
rect 15669 18717 15703 18751
rect 18705 18717 18739 18751
rect 20545 18717 20579 18751
rect 28549 18717 28583 18751
rect 21925 18649 21959 18683
rect 5917 18581 5951 18615
rect 7481 18581 7515 18615
rect 12725 18581 12759 18615
rect 14841 18581 14875 18615
rect 18981 18581 19015 18615
rect 25789 18581 25823 18615
rect 28825 18581 28859 18615
rect 1593 18377 1627 18411
rect 3525 18377 3559 18411
rect 10701 18377 10735 18411
rect 16681 18377 16715 18411
rect 21189 18377 21223 18411
rect 28365 18377 28399 18411
rect 28733 18377 28767 18411
rect 10425 18309 10459 18343
rect 17785 18309 17819 18343
rect 21465 18309 21499 18343
rect 1869 18241 1903 18275
rect 3801 18241 3835 18275
rect 6653 18241 6687 18275
rect 8125 18241 8159 18275
rect 9321 18241 9355 18275
rect 10149 18241 10183 18275
rect 13645 18241 13679 18275
rect 15485 18241 15519 18275
rect 17233 18241 17267 18275
rect 19901 18241 19935 18275
rect 22017 18241 22051 18275
rect 25513 18241 25547 18275
rect 29929 18241 29963 18275
rect 1685 18173 1719 18207
rect 1961 18173 1995 18207
rect 2053 18173 2087 18207
rect 2145 18173 2179 18207
rect 2329 18173 2363 18207
rect 2421 18173 2455 18207
rect 2605 18173 2639 18207
rect 3617 18173 3651 18207
rect 3893 18173 3927 18207
rect 3985 18173 4019 18207
rect 4077 18173 4111 18207
rect 4261 18173 4295 18207
rect 5917 18173 5951 18207
rect 6101 18173 6135 18207
rect 6193 18173 6227 18207
rect 6377 18173 6411 18207
rect 6469 18173 6503 18207
rect 6561 18173 6595 18207
rect 7665 18173 7699 18207
rect 7849 18173 7883 18207
rect 7941 18173 7975 18207
rect 8033 18173 8067 18207
rect 9413 18173 9447 18207
rect 9505 18173 9539 18207
rect 9965 18173 9999 18207
rect 10057 18173 10091 18207
rect 10333 18173 10367 18207
rect 10609 18173 10643 18207
rect 12725 18173 12759 18207
rect 13001 18173 13035 18207
rect 13185 18173 13219 18207
rect 13277 18173 13311 18207
rect 13553 18173 13587 18207
rect 14749 18173 14783 18207
rect 15025 18173 15059 18207
rect 15209 18173 15243 18207
rect 15301 18173 15335 18207
rect 15393 18173 15427 18207
rect 16773 18173 16807 18207
rect 16957 18173 16991 18207
rect 17049 18173 17083 18207
rect 17325 18173 17359 18207
rect 17417 18173 17451 18207
rect 17509 18173 17543 18207
rect 17693 18173 17727 18207
rect 18889 18173 18923 18207
rect 19441 18173 19475 18207
rect 19533 18173 19567 18207
rect 19625 18173 19659 18207
rect 19809 18173 19843 18207
rect 20085 18173 20119 18207
rect 21281 18173 21315 18207
rect 21557 18173 21591 18207
rect 21833 18173 21867 18207
rect 21925 18173 21959 18207
rect 22201 18173 22235 18207
rect 24501 18173 24535 18207
rect 24685 18173 24719 18207
rect 24777 18173 24811 18207
rect 25605 18173 25639 18207
rect 25973 18173 26007 18207
rect 26065 18173 26099 18207
rect 28457 18173 28491 18207
rect 28825 18173 28859 18207
rect 29101 18173 29135 18207
rect 29193 18173 29227 18207
rect 29377 18173 29411 18207
rect 29469 18173 29503 18207
rect 29745 18173 29779 18207
rect 29837 18173 29871 18207
rect 2697 18105 2731 18139
rect 4353 18105 4387 18139
rect 9873 18105 9907 18139
rect 12633 18105 12667 18139
rect 14657 18105 14691 18139
rect 19349 18105 19383 18139
rect 21741 18105 21775 18139
rect 26157 18105 26191 18139
rect 29653 18105 29687 18139
rect 5825 18037 5859 18071
rect 7573 18037 7607 18071
rect 9597 18037 9631 18071
rect 12909 18037 12943 18071
rect 14933 18037 14967 18071
rect 18981 18037 19015 18071
rect 20177 18037 20211 18071
rect 22293 18037 22327 18071
rect 24409 18037 24443 18071
rect 25881 18037 25915 18071
rect 2605 17833 2639 17867
rect 3893 17833 3927 17867
rect 9689 17833 9723 17867
rect 18061 17833 18095 17867
rect 19073 17833 19107 17867
rect 22293 17833 22327 17867
rect 25329 17833 25363 17867
rect 30021 17833 30055 17867
rect 4721 17765 4755 17799
rect 5549 17765 5583 17799
rect 7113 17765 7147 17799
rect 12817 17765 12851 17799
rect 13645 17765 13679 17799
rect 14841 17765 14875 17799
rect 20637 17765 20671 17799
rect 22569 17765 22603 17799
rect 25053 17765 25087 17799
rect 26801 17765 26835 17799
rect 1869 17697 1903 17731
rect 1961 17697 1995 17731
rect 2053 17697 2087 17731
rect 2237 17697 2271 17731
rect 2329 17697 2363 17731
rect 2513 17697 2547 17731
rect 3985 17697 4019 17731
rect 4077 17697 4111 17731
rect 4169 17697 4203 17731
rect 4353 17697 4387 17731
rect 4445 17697 4479 17731
rect 4629 17697 4663 17731
rect 5641 17697 5675 17731
rect 5825 17697 5859 17731
rect 5917 17697 5951 17731
rect 6101 17697 6135 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 6469 17697 6503 17731
rect 6745 17697 6779 17731
rect 6837 17697 6871 17731
rect 7021 17697 7055 17731
rect 7481 17697 7515 17731
rect 7573 17697 7607 17731
rect 7665 17697 7699 17731
rect 7941 17697 7975 17731
rect 8033 17697 8067 17731
rect 8217 17697 8251 17731
rect 8309 17697 8343 17731
rect 8493 17697 8527 17731
rect 8585 17697 8619 17731
rect 8769 17697 8803 17731
rect 8861 17697 8895 17731
rect 9045 17697 9079 17731
rect 9321 17697 9355 17731
rect 9597 17697 9631 17731
rect 12633 17697 12667 17731
rect 12909 17697 12943 17731
rect 13001 17697 13035 17731
rect 13461 17697 13495 17731
rect 13553 17697 13587 17731
rect 14933 17697 14967 17731
rect 15209 17697 15243 17731
rect 15393 17697 15427 17731
rect 15485 17697 15519 17731
rect 15577 17697 15611 17731
rect 17601 17697 17635 17731
rect 17693 17697 17727 17731
rect 17785 17697 17819 17731
rect 17969 17697 18003 17731
rect 18981 17697 19015 17731
rect 19625 17697 19659 17731
rect 19717 17697 19751 17731
rect 19809 17697 19843 17731
rect 19993 17697 20027 17731
rect 20453 17697 20487 17731
rect 20545 17697 20579 17731
rect 22109 17697 22143 17731
rect 22201 17697 22235 17731
rect 22661 17697 22695 17731
rect 22845 17697 22879 17731
rect 22937 17697 22971 17731
rect 23121 17697 23155 17731
rect 23213 17697 23247 17731
rect 23397 17697 23431 17731
rect 23489 17697 23523 17731
rect 23581 17697 23615 17731
rect 24041 17697 24075 17731
rect 24225 17697 24259 17731
rect 24317 17697 24351 17731
rect 24501 17697 24535 17731
rect 24593 17697 24627 17731
rect 24777 17697 24811 17731
rect 24869 17697 24903 17731
rect 24961 17697 24995 17731
rect 25237 17697 25271 17731
rect 25789 17697 25823 17731
rect 26249 17697 26283 17731
rect 26433 17697 26467 17731
rect 26525 17697 26559 17731
rect 26709 17697 26743 17731
rect 28089 17697 28123 17731
rect 29561 17697 29595 17731
rect 29653 17697 29687 17731
rect 29745 17697 29779 17731
rect 29929 17697 29963 17731
rect 9137 17629 9171 17663
rect 13369 17629 13403 17663
rect 15669 17629 15703 17663
rect 17509 17629 17543 17663
rect 19533 17629 19567 17663
rect 20085 17629 20119 17663
rect 22017 17629 22051 17663
rect 23673 17629 23707 17663
rect 25881 17629 25915 17663
rect 29469 17629 29503 17663
rect 13093 17561 13127 17595
rect 1777 17493 1811 17527
rect 7389 17493 7423 17527
rect 9413 17493 9447 17527
rect 12541 17493 12575 17527
rect 15117 17493 15151 17527
rect 20361 17493 20395 17527
rect 23949 17493 23983 17527
rect 26157 17493 26191 17527
rect 28181 17493 28215 17527
rect 1225 17289 1259 17323
rect 3985 17289 4019 17323
rect 9045 17289 9079 17323
rect 17601 17289 17635 17323
rect 22937 17289 22971 17323
rect 24869 17289 24903 17323
rect 30205 17289 30239 17323
rect 4813 17153 4847 17187
rect 7849 17153 7883 17187
rect 12633 17153 12667 17187
rect 14841 17153 14875 17187
rect 20361 17153 20395 17187
rect 1317 17085 1351 17119
rect 1593 17085 1627 17119
rect 1777 17085 1811 17119
rect 1869 17085 1903 17119
rect 2053 17085 2087 17119
rect 2145 17085 2179 17119
rect 2329 17085 2363 17119
rect 2421 17085 2455 17119
rect 2605 17085 2639 17119
rect 2697 17085 2731 17119
rect 2881 17085 2915 17119
rect 2973 17085 3007 17119
rect 3341 17085 3375 17119
rect 3433 17085 3467 17119
rect 3709 17085 3743 17119
rect 3801 17085 3835 17119
rect 4077 17085 4111 17119
rect 4261 17085 4295 17119
rect 4353 17085 4387 17119
rect 4629 17085 4663 17119
rect 4905 17085 4939 17119
rect 5181 17085 5215 17119
rect 7665 17085 7699 17119
rect 7757 17085 7791 17119
rect 9137 17085 9171 17119
rect 9321 17085 9355 17119
rect 9413 17085 9447 17119
rect 9689 17085 9723 17119
rect 9873 17085 9907 17119
rect 9965 17085 9999 17119
rect 10149 17085 10183 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 10793 17085 10827 17119
rect 11069 17085 11103 17119
rect 11253 17085 11287 17119
rect 11345 17085 11379 17119
rect 11529 17085 11563 17119
rect 11621 17085 11655 17119
rect 11805 17085 11839 17119
rect 11897 17085 11931 17119
rect 12081 17085 12115 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 12541 17085 12575 17119
rect 13829 17085 13863 17119
rect 13921 17085 13955 17119
rect 14105 17085 14139 17119
rect 14197 17085 14231 17119
rect 14473 17085 14507 17119
rect 14565 17085 14599 17119
rect 14749 17085 14783 17119
rect 15025 17085 15059 17119
rect 15301 17085 15335 17119
rect 15393 17085 15427 17119
rect 15761 17085 15795 17119
rect 15853 17085 15887 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 16313 17085 16347 17119
rect 16405 17085 16439 17119
rect 16589 17085 16623 17119
rect 17693 17085 17727 17119
rect 17877 17085 17911 17119
rect 17969 17085 18003 17119
rect 18153 17085 18187 17119
rect 18245 17085 18279 17119
rect 18429 17085 18463 17119
rect 18521 17085 18555 17119
rect 18797 17085 18831 17119
rect 18889 17085 18923 17119
rect 19073 17085 19107 17119
rect 19165 17085 19199 17119
rect 19257 17085 19291 17119
rect 20269 17085 20303 17119
rect 20729 17085 20763 17119
rect 20821 17085 20855 17119
rect 20913 17085 20947 17119
rect 21097 17085 21131 17119
rect 23029 17085 23063 17119
rect 24225 17085 24259 17119
rect 24317 17085 24351 17119
rect 24501 17085 24535 17119
rect 24593 17085 24627 17119
rect 24777 17085 24811 17119
rect 26341 17085 26375 17119
rect 26433 17085 26467 17119
rect 26617 17085 26651 17119
rect 26709 17085 26743 17119
rect 26893 17085 26927 17119
rect 26985 17085 27019 17119
rect 27169 17085 27203 17119
rect 27261 17085 27295 17119
rect 27445 17085 27479 17119
rect 27537 17085 27571 17119
rect 27721 17085 27755 17119
rect 27813 17085 27847 17119
rect 27997 17085 28031 17119
rect 28089 17085 28123 17119
rect 28273 17085 28307 17119
rect 28365 17085 28399 17119
rect 28549 17085 28583 17119
rect 29009 17085 29043 17119
rect 29101 17085 29135 17119
rect 29285 17085 29319 17119
rect 29377 17085 29411 17119
rect 29561 17085 29595 17119
rect 29653 17085 29687 17119
rect 29837 17085 29871 17119
rect 30113 17085 30147 17119
rect 4537 17017 4571 17051
rect 5089 17017 5123 17051
rect 12357 17017 12391 17051
rect 19349 17017 19383 17051
rect 21189 17017 21223 17051
rect 1501 16949 1535 16983
rect 7573 16949 7607 16983
rect 9597 16949 9631 16983
rect 10977 16949 11011 16983
rect 15117 16949 15151 16983
rect 16681 16949 16715 16983
rect 20637 16949 20671 16983
rect 28641 16949 28675 16983
rect 29929 16949 29963 16983
rect 1869 16745 1903 16779
rect 4905 16745 4939 16779
rect 5273 16745 5307 16779
rect 9873 16745 9907 16779
rect 11253 16745 11287 16779
rect 13645 16745 13679 16779
rect 18797 16745 18831 16779
rect 24501 16745 24535 16779
rect 27997 16745 28031 16779
rect 29285 16745 29319 16779
rect 6469 16677 6503 16711
rect 8217 16677 8251 16711
rect 10149 16677 10183 16711
rect 14197 16677 14231 16711
rect 15485 16677 15519 16711
rect 17325 16677 17359 16711
rect 19625 16677 19659 16711
rect 24225 16677 24259 16711
rect 25053 16677 25087 16711
rect 29837 16677 29871 16711
rect 1777 16609 1811 16643
rect 4261 16609 4295 16643
rect 4353 16609 4387 16643
rect 4537 16609 4571 16643
rect 4629 16609 4663 16643
rect 4813 16609 4847 16643
rect 5365 16609 5399 16643
rect 5549 16609 5583 16643
rect 5641 16609 5675 16643
rect 5917 16609 5951 16643
rect 6009 16609 6043 16643
rect 6101 16609 6135 16643
rect 6193 16609 6227 16643
rect 6377 16609 6411 16643
rect 7757 16609 7791 16643
rect 7941 16609 7975 16643
rect 8033 16609 8067 16643
rect 8125 16609 8159 16643
rect 9321 16609 9355 16643
rect 9505 16609 9539 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 10057 16609 10091 16643
rect 11161 16609 11195 16643
rect 13185 16609 13219 16643
rect 13277 16609 13311 16643
rect 13737 16609 13771 16643
rect 13921 16609 13955 16643
rect 14013 16609 14047 16643
rect 14105 16609 14139 16643
rect 15301 16609 15335 16643
rect 15393 16609 15427 16643
rect 16681 16609 16715 16643
rect 16773 16609 16807 16643
rect 17141 16609 17175 16643
rect 17233 16609 17267 16643
rect 18889 16609 18923 16643
rect 18981 16609 19015 16643
rect 19073 16609 19107 16643
rect 19257 16609 19291 16643
rect 19349 16609 19383 16643
rect 19533 16609 19567 16643
rect 20729 16609 20763 16643
rect 20821 16609 20855 16643
rect 21281 16609 21315 16643
rect 21373 16609 21407 16643
rect 21557 16609 21591 16643
rect 21649 16609 21683 16643
rect 21833 16609 21867 16643
rect 21925 16609 21959 16643
rect 22109 16609 22143 16643
rect 22201 16609 22235 16643
rect 22385 16609 22419 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 24041 16609 24075 16643
rect 24317 16609 24351 16643
rect 24409 16609 24443 16643
rect 24777 16609 24811 16643
rect 24869 16609 24903 16643
rect 24961 16609 24995 16643
rect 25513 16609 25547 16643
rect 25697 16609 25731 16643
rect 25789 16609 25823 16643
rect 25973 16609 26007 16643
rect 26065 16609 26099 16643
rect 28089 16609 28123 16643
rect 29377 16609 29411 16643
rect 29929 16609 29963 16643
rect 7665 16405 7699 16439
rect 9229 16405 9263 16439
rect 15209 16405 15243 16439
rect 17049 16405 17083 16439
rect 22753 16405 22787 16439
rect 23949 16405 23983 16439
rect 25421 16405 25455 16439
rect 3893 16201 3927 16235
rect 6193 16201 6227 16235
rect 12817 16201 12851 16235
rect 18889 16201 18923 16235
rect 24225 16201 24259 16235
rect 24777 16201 24811 16235
rect 25973 16201 26007 16235
rect 30205 16201 30239 16235
rect 6469 16065 6503 16099
rect 7297 16065 7331 16099
rect 9689 16065 9723 16099
rect 11161 16065 11195 16099
rect 13921 16065 13955 16099
rect 15945 16065 15979 16099
rect 17693 16065 17727 16099
rect 19165 16065 19199 16099
rect 22109 16065 22143 16099
rect 3985 15997 4019 16031
rect 4261 15997 4295 16031
rect 4445 15997 4479 16031
rect 4537 15997 4571 16031
rect 4629 15997 4663 16031
rect 4721 15997 4755 16031
rect 4905 15997 4939 16031
rect 6285 15997 6319 16031
rect 6561 15997 6595 16031
rect 6653 15997 6687 16031
rect 6745 15997 6779 16031
rect 6929 15997 6963 16031
rect 7389 15997 7423 16031
rect 7481 15997 7515 16031
rect 7573 15997 7607 16031
rect 7757 15997 7791 16031
rect 7849 15997 7883 16031
rect 8033 15997 8067 16031
rect 8125 15997 8159 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 8677 15997 8711 16031
rect 9229 15997 9263 16031
rect 9321 15997 9355 16031
rect 9597 15997 9631 16031
rect 11069 15997 11103 16031
rect 11621 15997 11655 16031
rect 11713 15997 11747 16031
rect 12909 15997 12943 16031
rect 13185 15997 13219 16031
rect 13553 15997 13587 16031
rect 13645 15997 13679 16031
rect 13829 15997 13863 16031
rect 14933 15997 14967 16031
rect 15209 15997 15243 16031
rect 15393 15997 15427 16031
rect 15485 15997 15519 16031
rect 15669 15997 15703 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 16957 15997 16991 16031
rect 17233 15997 17267 16031
rect 17417 15997 17451 16031
rect 17509 15997 17543 16031
rect 17601 15997 17635 16031
rect 18981 15997 19015 16031
rect 19257 15997 19291 16031
rect 19349 15997 19383 16031
rect 19441 15997 19475 16031
rect 19625 15997 19659 16031
rect 22201 15997 22235 16031
rect 22293 15997 22327 16031
rect 22385 15997 22419 16031
rect 22569 15997 22603 16031
rect 22661 15997 22695 16031
rect 22845 15997 22879 16031
rect 22937 15997 22971 16031
rect 23121 15997 23155 16031
rect 23213 15997 23247 16031
rect 23397 15997 23431 16031
rect 24133 15997 24167 16031
rect 24869 15997 24903 16031
rect 25053 15997 25087 16031
rect 25145 15997 25179 16031
rect 25329 15997 25363 16031
rect 25421 15997 25455 16031
rect 26065 15997 26099 16031
rect 26249 15997 26283 16031
rect 26341 15997 26375 16031
rect 26525 15997 26559 16031
rect 26617 15997 26651 16031
rect 26801 15997 26835 16031
rect 26893 15997 26927 16031
rect 27077 15997 27111 16031
rect 27169 15997 27203 16031
rect 27353 15997 27387 16031
rect 27445 15997 27479 16031
rect 27629 15997 27663 16031
rect 27721 15997 27755 16031
rect 27905 15997 27939 16031
rect 27997 15997 28031 16031
rect 28181 15997 28215 16031
rect 28273 15997 28307 16031
rect 28457 15997 28491 16031
rect 28549 15997 28583 16031
rect 28733 15997 28767 16031
rect 28825 15997 28859 16031
rect 29101 15997 29135 16031
rect 29193 15997 29227 16031
rect 29377 15997 29411 16031
rect 29469 15997 29503 16031
rect 29653 15997 29687 16031
rect 29745 15997 29779 16031
rect 29929 15997 29963 16031
rect 30021 15997 30055 16031
rect 30113 15997 30147 16031
rect 30389 15997 30423 16031
rect 4169 15929 4203 15963
rect 7021 15929 7055 15963
rect 8769 15929 8803 15963
rect 11805 15929 11839 15963
rect 13093 15929 13127 15963
rect 14841 15929 14875 15963
rect 16865 15929 16899 15963
rect 19717 15929 19751 15963
rect 30481 15929 30515 15963
rect 4997 15861 5031 15895
rect 9137 15861 9171 15895
rect 9413 15861 9447 15895
rect 11529 15861 11563 15895
rect 15117 15861 15151 15895
rect 17141 15861 17175 15895
rect 23489 15861 23523 15895
rect 4905 15657 4939 15691
rect 6929 15657 6963 15691
rect 11069 15657 11103 15691
rect 13185 15657 13219 15691
rect 19809 15657 19843 15691
rect 30113 15657 30147 15691
rect 11345 15589 11379 15623
rect 12909 15589 12943 15623
rect 23581 15589 23615 15623
rect 29285 15589 29319 15623
rect 3985 15521 4019 15555
rect 4077 15521 4111 15555
rect 4261 15521 4295 15555
rect 4353 15521 4387 15555
rect 4537 15521 4571 15555
rect 4629 15521 4663 15555
rect 4813 15521 4847 15555
rect 6285 15521 6319 15555
rect 6377 15521 6411 15555
rect 6561 15521 6595 15555
rect 6653 15521 6687 15555
rect 6837 15521 6871 15555
rect 8953 15521 8987 15555
rect 9045 15521 9079 15555
rect 9413 15521 9447 15555
rect 9505 15521 9539 15555
rect 9781 15521 9815 15555
rect 9873 15521 9907 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 10333 15521 10367 15555
rect 10425 15521 10459 15555
rect 10609 15521 10643 15555
rect 11161 15521 11195 15555
rect 11253 15521 11287 15555
rect 11621 15521 11655 15555
rect 11713 15521 11747 15555
rect 11897 15521 11931 15555
rect 11989 15521 12023 15555
rect 12173 15521 12207 15555
rect 12265 15521 12299 15555
rect 12449 15521 12483 15555
rect 13001 15521 13035 15555
rect 13093 15521 13127 15555
rect 13369 15521 13403 15555
rect 14841 15521 14875 15555
rect 15025 15521 15059 15555
rect 15117 15521 15151 15555
rect 15301 15521 15335 15555
rect 15393 15521 15427 15555
rect 15577 15521 15611 15555
rect 15669 15521 15703 15555
rect 15761 15521 15795 15555
rect 16957 15521 16991 15555
rect 17141 15521 17175 15555
rect 17233 15521 17267 15555
rect 17417 15521 17451 15555
rect 17509 15521 17543 15555
rect 17601 15521 17635 15555
rect 19073 15521 19107 15555
rect 19165 15521 19199 15555
rect 19257 15521 19291 15555
rect 19441 15521 19475 15555
rect 19533 15521 19567 15555
rect 19717 15521 19751 15555
rect 22109 15521 22143 15555
rect 23121 15521 23155 15555
rect 23213 15521 23247 15555
rect 23305 15521 23339 15555
rect 23489 15521 23523 15555
rect 23949 15521 23983 15555
rect 24041 15521 24075 15555
rect 24317 15521 24351 15555
rect 29377 15521 29411 15555
rect 29469 15521 29503 15555
rect 29561 15521 29595 15555
rect 29745 15521 29779 15555
rect 29837 15521 29871 15555
rect 30021 15521 30055 15555
rect 8861 15453 8895 15487
rect 10701 15453 10735 15487
rect 13461 15453 13495 15487
rect 15853 15453 15887 15487
rect 17693 15453 17727 15487
rect 18981 15453 19015 15487
rect 23029 15453 23063 15487
rect 24133 15453 24167 15487
rect 12541 15385 12575 15419
rect 23857 15385 23891 15419
rect 9137 15317 9171 15351
rect 14749 15317 14783 15351
rect 16865 15317 16899 15351
rect 22201 15317 22235 15351
rect 24409 15317 24443 15351
rect 3801 15113 3835 15147
rect 6009 15113 6043 15147
rect 19625 15113 19659 15147
rect 29929 15113 29963 15147
rect 4353 14977 4387 15011
rect 6745 14977 6779 15011
rect 7573 14977 7607 15011
rect 9413 14977 9447 15011
rect 14933 14977 14967 15011
rect 17325 14977 17359 15011
rect 18429 14977 18463 15011
rect 22845 14977 22879 15011
rect 23305 14977 23339 15011
rect 2329 14909 2363 14943
rect 2513 14909 2547 14943
rect 2605 14909 2639 14943
rect 2789 14909 2823 14943
rect 2881 14909 2915 14943
rect 3341 14909 3375 14943
rect 3433 14909 3467 14943
rect 3893 14909 3927 14943
rect 4077 14909 4111 14943
rect 4169 14909 4203 14943
rect 4445 14909 4479 14943
rect 4629 14909 4663 14943
rect 4721 14909 4755 14943
rect 4905 14909 4939 14943
rect 4997 14909 5031 14943
rect 5181 14909 5215 14943
rect 5273 14909 5307 14943
rect 5457 14909 5491 14943
rect 5549 14909 5583 14943
rect 5733 14909 5767 14943
rect 5825 14909 5859 14943
rect 6101 14909 6135 14943
rect 6285 14909 6319 14943
rect 6377 14909 6411 14943
rect 6837 14909 6871 14943
rect 7113 14909 7147 14943
rect 7205 14909 7239 14943
rect 7665 14909 7699 14943
rect 7757 14909 7791 14943
rect 9229 14909 9263 14943
rect 9321 14909 9355 14943
rect 10701 14909 10735 14943
rect 11713 14909 11747 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 14749 14909 14783 14943
rect 14841 14909 14875 14943
rect 16589 14909 16623 14943
rect 16773 14909 16807 14943
rect 16865 14909 16899 14943
rect 17049 14909 17083 14943
rect 17141 14909 17175 14943
rect 17233 14909 17267 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 18797 14909 18831 14943
rect 18981 14909 19015 14943
rect 19073 14909 19107 14943
rect 19257 14909 19291 14943
rect 19349 14909 19383 14943
rect 19533 14909 19567 14943
rect 20453 14909 20487 14943
rect 20637 14909 20671 14943
rect 20729 14909 20763 14943
rect 20913 14909 20947 14943
rect 21005 14909 21039 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 21465 14909 21499 14943
rect 21557 14909 21591 14943
rect 21741 14909 21775 14943
rect 21833 14909 21867 14943
rect 22017 14909 22051 14943
rect 22109 14909 22143 14943
rect 22293 14909 22327 14943
rect 22385 14909 22419 14943
rect 22569 14909 22603 14943
rect 22661 14909 22695 14943
rect 22753 14909 22787 14943
rect 23397 14909 23431 14943
rect 23581 14909 23615 14943
rect 23673 14909 23707 14943
rect 24225 14909 24259 14943
rect 24317 14909 24351 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 29009 14909 29043 14943
rect 29101 14909 29135 14943
rect 29285 14909 29319 14943
rect 29377 14909 29411 14943
rect 29561 14909 29595 14943
rect 29653 14909 29687 14943
rect 29837 14909 29871 14943
rect 30573 14909 30607 14943
rect 7849 14841 7883 14875
rect 24685 14841 24719 14875
rect 2237 14773 2271 14807
rect 9137 14773 9171 14807
rect 10793 14773 10827 14807
rect 11805 14773 11839 14807
rect 14381 14773 14415 14807
rect 16497 14773 16531 14807
rect 20361 14773 20395 14807
rect 24133 14773 24167 14807
rect 30481 14773 30515 14807
rect 2881 14569 2915 14603
rect 4353 14569 4387 14603
rect 6469 14569 6503 14603
rect 7665 14569 7699 14603
rect 10425 14569 10459 14603
rect 11529 14569 11563 14603
rect 18613 14569 18647 14603
rect 22109 14569 22143 14603
rect 29101 14569 29135 14603
rect 31033 14569 31067 14603
rect 2605 14501 2639 14535
rect 9045 14501 9079 14535
rect 14841 14501 14875 14535
rect 16313 14501 16347 14535
rect 22937 14501 22971 14535
rect 1869 14433 1903 14467
rect 2145 14433 2179 14467
rect 2329 14433 2363 14467
rect 2421 14433 2455 14467
rect 2513 14433 2547 14467
rect 2789 14433 2823 14467
rect 4169 14433 4203 14467
rect 4261 14433 4295 14467
rect 6101 14433 6135 14467
rect 6193 14433 6227 14467
rect 6377 14433 6411 14467
rect 7757 14433 7791 14467
rect 7941 14433 7975 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 8309 14433 8343 14467
rect 8493 14433 8527 14467
rect 8585 14433 8619 14467
rect 8769 14433 8803 14467
rect 8861 14433 8895 14467
rect 9137 14433 9171 14467
rect 9229 14433 9263 14467
rect 9505 14433 9539 14467
rect 10517 14433 10551 14467
rect 10701 14433 10735 14467
rect 10793 14433 10827 14467
rect 11345 14433 11379 14467
rect 11621 14433 11655 14467
rect 11805 14433 11839 14467
rect 11897 14433 11931 14467
rect 12081 14433 12115 14467
rect 12173 14433 12207 14467
rect 12357 14433 12391 14467
rect 12449 14433 12483 14467
rect 12633 14433 12667 14467
rect 12725 14433 12759 14467
rect 12909 14433 12943 14467
rect 13001 14433 13035 14467
rect 13185 14433 13219 14467
rect 13277 14433 13311 14467
rect 13461 14433 13495 14467
rect 13553 14433 13587 14467
rect 13737 14433 13771 14467
rect 13829 14433 13863 14467
rect 14013 14433 14047 14467
rect 14105 14433 14139 14467
rect 14381 14433 14415 14467
rect 14473 14433 14507 14467
rect 14565 14433 14599 14467
rect 14749 14433 14783 14467
rect 15393 14433 15427 14467
rect 15577 14433 15611 14467
rect 15669 14433 15703 14467
rect 15853 14433 15887 14467
rect 15945 14433 15979 14467
rect 16405 14433 16439 14467
rect 16497 14433 16531 14467
rect 17601 14433 17635 14467
rect 17693 14433 17727 14467
rect 17785 14433 17819 14467
rect 17969 14433 18003 14467
rect 18061 14433 18095 14467
rect 18245 14433 18279 14467
rect 18337 14433 18371 14467
rect 18521 14433 18555 14467
rect 20453 14433 20487 14467
rect 20637 14433 20671 14467
rect 20729 14433 20763 14467
rect 20821 14433 20855 14467
rect 22201 14433 22235 14467
rect 22477 14433 22511 14467
rect 22569 14433 22603 14467
rect 22661 14433 22695 14467
rect 22845 14433 22879 14467
rect 24133 14433 24167 14467
rect 24225 14433 24259 14467
rect 24317 14433 24351 14467
rect 24501 14433 24535 14467
rect 24593 14433 24627 14467
rect 24777 14433 24811 14467
rect 24869 14433 24903 14467
rect 25053 14433 25087 14467
rect 29193 14433 29227 14467
rect 29377 14433 29411 14467
rect 29469 14433 29503 14467
rect 29653 14433 29687 14467
rect 29745 14433 29779 14467
rect 29929 14433 29963 14467
rect 30021 14433 30055 14467
rect 30205 14433 30239 14467
rect 30297 14433 30331 14467
rect 30389 14433 30423 14467
rect 30849 14433 30883 14467
rect 30941 14433 30975 14467
rect 1777 14365 1811 14399
rect 4077 14365 4111 14399
rect 9321 14365 9355 14399
rect 14289 14365 14323 14399
rect 16589 14365 16623 14399
rect 17509 14365 17543 14399
rect 20913 14365 20947 14399
rect 22385 14365 22419 14399
rect 24041 14365 24075 14399
rect 30481 14365 30515 14399
rect 30757 14365 30791 14399
rect 9597 14297 9631 14331
rect 2053 14229 2087 14263
rect 11253 14229 11287 14263
rect 15301 14229 15335 14263
rect 20361 14229 20395 14263
rect 25145 14229 25179 14263
rect 4905 14025 4939 14059
rect 11345 14025 11379 14059
rect 17785 14025 17819 14059
rect 23213 14025 23247 14059
rect 31125 14025 31159 14059
rect 19165 13957 19199 13991
rect 2605 13889 2639 13923
rect 7021 13889 7055 13923
rect 16313 13889 16347 13923
rect 17233 13889 17267 13923
rect 21097 13889 21131 13923
rect 22109 13889 22143 13923
rect 25053 13889 25087 13923
rect 30573 13889 30607 13923
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 2421 13821 2455 13855
rect 2513 13821 2547 13855
rect 3985 13821 4019 13855
rect 4077 13821 4111 13855
rect 4261 13821 4295 13855
rect 4353 13821 4387 13855
rect 4537 13821 4571 13855
rect 4629 13821 4663 13855
rect 4813 13821 4847 13855
rect 5917 13821 5951 13855
rect 6101 13821 6135 13855
rect 6193 13821 6227 13855
rect 6377 13821 6411 13855
rect 6469 13821 6503 13855
rect 6653 13821 6687 13855
rect 6745 13821 6779 13855
rect 6929 13821 6963 13855
rect 10609 13821 10643 13855
rect 10793 13821 10827 13855
rect 10885 13821 10919 13855
rect 11253 13821 11287 13855
rect 11805 13821 11839 13855
rect 15577 13821 15611 13855
rect 15761 13821 15795 13855
rect 15853 13821 15887 13855
rect 16037 13821 16071 13855
rect 16129 13821 16163 13855
rect 16221 13821 16255 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 17509 13821 17543 13855
rect 17693 13821 17727 13855
rect 19257 13821 19291 13855
rect 19441 13821 19475 13855
rect 19533 13821 19567 13855
rect 19717 13821 19751 13855
rect 19809 13821 19843 13855
rect 19993 13821 20027 13855
rect 20085 13821 20119 13855
rect 20269 13821 20303 13855
rect 20361 13821 20395 13855
rect 20545 13821 20579 13855
rect 20637 13821 20671 13855
rect 20821 13821 20855 13855
rect 20913 13821 20947 13855
rect 21005 13821 21039 13855
rect 22201 13821 22235 13855
rect 22293 13821 22327 13855
rect 22385 13821 22419 13855
rect 22569 13821 22603 13855
rect 22661 13821 22695 13855
rect 22845 13821 22879 13855
rect 22937 13821 22971 13855
rect 23121 13821 23155 13855
rect 25145 13821 25179 13855
rect 25237 13821 25271 13855
rect 25329 13821 25363 13855
rect 25513 13821 25547 13855
rect 25605 13821 25639 13855
rect 25789 13821 25823 13855
rect 25881 13821 25915 13855
rect 26065 13821 26099 13855
rect 26157 13821 26191 13855
rect 26341 13821 26375 13855
rect 26433 13821 26467 13855
rect 26617 13821 26651 13855
rect 26709 13821 26743 13855
rect 26893 13821 26927 13855
rect 26985 13821 27019 13855
rect 27169 13821 27203 13855
rect 27261 13821 27295 13855
rect 27445 13821 27479 13855
rect 27537 13821 27571 13855
rect 27721 13821 27755 13855
rect 27813 13821 27847 13855
rect 27997 13821 28031 13855
rect 28089 13821 28123 13855
rect 28273 13821 28307 13855
rect 28365 13821 28399 13855
rect 28549 13821 28583 13855
rect 28641 13821 28675 13855
rect 29009 13821 29043 13855
rect 30665 13821 30699 13855
rect 30757 13821 30791 13855
rect 30849 13821 30883 13855
rect 31033 13821 31067 13855
rect 2053 13685 2087 13719
rect 5825 13685 5859 13719
rect 10517 13685 10551 13719
rect 11897 13685 11931 13719
rect 15485 13685 15519 13719
rect 29101 13685 29135 13719
rect 4077 13481 4111 13515
rect 6193 13481 6227 13515
rect 6653 13481 6687 13515
rect 11805 13481 11839 13515
rect 17877 13481 17911 13515
rect 20361 13481 20395 13515
rect 22753 13481 22787 13515
rect 31217 13481 31251 13515
rect 1869 13413 1903 13447
rect 2973 13413 3007 13447
rect 4905 13413 4939 13447
rect 13001 13413 13035 13447
rect 15209 13413 15243 13447
rect 18153 13413 18187 13447
rect 1961 13345 1995 13379
rect 2053 13345 2087 13379
rect 2513 13345 2547 13379
rect 2697 13345 2731 13379
rect 2789 13345 2823 13379
rect 2881 13345 2915 13379
rect 4169 13345 4203 13379
rect 4261 13345 4295 13379
rect 4353 13345 4387 13379
rect 4537 13345 4571 13379
rect 4629 13345 4663 13379
rect 4813 13345 4847 13379
rect 6101 13345 6135 13379
rect 6745 13345 6779 13379
rect 6929 13345 6963 13379
rect 7021 13345 7055 13379
rect 7297 13345 7331 13379
rect 7481 13345 7515 13379
rect 7573 13345 7607 13379
rect 7757 13345 7791 13379
rect 7849 13345 7883 13379
rect 8033 13345 8067 13379
rect 8125 13345 8159 13379
rect 8309 13345 8343 13379
rect 8401 13345 8435 13379
rect 8585 13345 8619 13379
rect 8677 13345 8711 13379
rect 8861 13345 8895 13379
rect 8953 13345 8987 13379
rect 9137 13345 9171 13379
rect 9229 13345 9263 13379
rect 9413 13345 9447 13379
rect 9505 13345 9539 13379
rect 9689 13345 9723 13379
rect 9781 13345 9815 13379
rect 9965 13345 9999 13379
rect 10057 13345 10091 13379
rect 10241 13345 10275 13379
rect 10333 13345 10367 13379
rect 10517 13345 10551 13379
rect 10609 13345 10643 13379
rect 10977 13345 11011 13379
rect 11621 13345 11655 13379
rect 11897 13345 11931 13379
rect 12081 13345 12115 13379
rect 12173 13345 12207 13379
rect 12357 13345 12391 13379
rect 12449 13345 12483 13379
rect 12633 13345 12667 13379
rect 12725 13345 12759 13379
rect 13093 13345 13127 13379
rect 13185 13345 13219 13379
rect 15301 13345 15335 13379
rect 15577 13345 15611 13379
rect 15761 13345 15795 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 17417 13345 17451 13379
rect 17509 13345 17543 13379
rect 17601 13345 17635 13379
rect 17785 13345 17819 13379
rect 18245 13345 18279 13379
rect 18429 13345 18463 13379
rect 18521 13345 18555 13379
rect 18705 13345 18739 13379
rect 18797 13345 18831 13379
rect 18981 13345 19015 13379
rect 19073 13345 19107 13379
rect 19257 13345 19291 13379
rect 19349 13345 19383 13379
rect 19441 13345 19475 13379
rect 20269 13345 20303 13379
rect 21557 13345 21591 13379
rect 21649 13345 21683 13379
rect 21833 13345 21867 13379
rect 21925 13345 21959 13379
rect 22109 13345 22143 13379
rect 22201 13345 22235 13379
rect 22385 13345 22419 13379
rect 22477 13345 22511 13379
rect 22661 13345 22695 13379
rect 25053 13345 25087 13379
rect 25237 13345 25271 13379
rect 25329 13345 25363 13379
rect 25605 13345 25639 13379
rect 25697 13345 25731 13379
rect 25881 13345 25915 13379
rect 25973 13345 26007 13379
rect 26617 13345 26651 13379
rect 28457 13345 28491 13379
rect 28641 13345 28675 13379
rect 28733 13345 28767 13379
rect 28917 13345 28951 13379
rect 29009 13345 29043 13379
rect 29101 13345 29135 13379
rect 30205 13345 30239 13379
rect 30297 13345 30331 13379
rect 30389 13345 30423 13379
rect 30573 13345 30607 13379
rect 30665 13345 30699 13379
rect 30849 13345 30883 13379
rect 30941 13345 30975 13379
rect 31125 13345 31159 13379
rect 2145 13277 2179 13311
rect 11069 13277 11103 13311
rect 13277 13277 13311 13311
rect 16221 13277 16255 13311
rect 17325 13277 17359 13311
rect 19533 13277 19567 13311
rect 29193 13277 29227 13311
rect 30113 13277 30147 13311
rect 2421 13141 2455 13175
rect 7205 13141 7239 13175
rect 11529 13141 11563 13175
rect 15485 13141 15519 13175
rect 24961 13141 24995 13175
rect 26525 13141 26559 13175
rect 28365 13141 28399 13175
rect 4169 12937 4203 12971
rect 7481 12937 7515 12971
rect 13921 12937 13955 12971
rect 21649 12937 21683 12971
rect 26157 12937 26191 12971
rect 26893 12937 26927 12971
rect 30757 12937 30791 12971
rect 2329 12801 2363 12835
rect 3341 12801 3375 12835
rect 5365 12801 5399 12835
rect 13277 12801 13311 12835
rect 15761 12801 15795 12835
rect 19073 12801 19107 12835
rect 22477 12801 22511 12835
rect 25421 12801 25455 12835
rect 26617 12801 26651 12835
rect 2421 12733 2455 12767
rect 2513 12733 2547 12767
rect 2973 12733 3007 12767
rect 3249 12733 3283 12767
rect 4261 12733 4295 12767
rect 4445 12733 4479 12767
rect 4537 12733 4571 12767
rect 4721 12733 4755 12767
rect 4813 12733 4847 12767
rect 4997 12733 5031 12767
rect 5089 12733 5123 12767
rect 5273 12733 5307 12767
rect 6193 12733 6227 12767
rect 7389 12733 7423 12767
rect 11621 12733 11655 12767
rect 11805 12733 11839 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 13645 12733 13679 12767
rect 13829 12733 13863 12767
rect 15301 12733 15335 12767
rect 15485 12733 15519 12767
rect 15577 12733 15611 12767
rect 15669 12733 15703 12767
rect 19165 12733 19199 12767
rect 19257 12733 19291 12767
rect 19349 12733 19383 12767
rect 19533 12733 19567 12767
rect 19625 12733 19659 12767
rect 19809 12733 19843 12767
rect 19901 12733 19935 12767
rect 20085 12733 20119 12767
rect 20177 12733 20211 12767
rect 20361 12733 20395 12767
rect 21741 12733 21775 12767
rect 21833 12733 21867 12767
rect 21925 12733 21959 12767
rect 22109 12733 22143 12767
rect 22201 12733 22235 12767
rect 22385 12733 22419 12767
rect 24409 12733 24443 12767
rect 24593 12733 24627 12767
rect 24685 12733 24719 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 25145 12733 25179 12767
rect 25237 12733 25271 12767
rect 25329 12733 25363 12767
rect 26249 12733 26283 12767
rect 26709 12733 26743 12767
rect 26801 12733 26835 12767
rect 27077 12733 27111 12767
rect 28365 12733 28399 12767
rect 28549 12733 28583 12767
rect 28641 12733 28675 12767
rect 29009 12733 29043 12767
rect 30021 12733 30055 12767
rect 30113 12733 30147 12767
rect 30205 12733 30239 12767
rect 30389 12733 30423 12767
rect 30481 12733 30515 12767
rect 30665 12733 30699 12767
rect 2605 12665 2639 12699
rect 12081 12665 12115 12699
rect 27169 12665 27203 12699
rect 29101 12665 29135 12699
rect 29929 12665 29963 12699
rect 2881 12597 2915 12631
rect 6101 12597 6135 12631
rect 11529 12597 11563 12631
rect 15209 12597 15243 12631
rect 20453 12597 20487 12631
rect 24317 12597 24351 12631
rect 28273 12597 28307 12631
rect 4997 12393 5031 12427
rect 13921 12393 13955 12427
rect 19625 12393 19659 12427
rect 21925 12393 21959 12427
rect 27077 12393 27111 12427
rect 30849 12393 30883 12427
rect 3709 12325 3743 12359
rect 9321 12325 9355 12359
rect 11989 12325 12023 12359
rect 14933 12325 14967 12359
rect 20177 12325 20211 12359
rect 22201 12325 22235 12359
rect 30573 12325 30607 12359
rect 2789 12257 2823 12291
rect 3249 12257 3283 12291
rect 3433 12257 3467 12291
rect 3525 12257 3559 12291
rect 3617 12257 3651 12291
rect 5089 12257 5123 12291
rect 5273 12257 5307 12291
rect 5365 12257 5399 12291
rect 5549 12257 5583 12291
rect 5641 12257 5675 12291
rect 6193 12257 6227 12291
rect 6377 12257 6411 12291
rect 6469 12257 6503 12291
rect 6653 12257 6687 12291
rect 6745 12257 6779 12291
rect 6929 12257 6963 12291
rect 7021 12257 7055 12291
rect 7205 12257 7239 12291
rect 7297 12257 7331 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 7757 12257 7791 12291
rect 7849 12257 7883 12291
rect 8033 12257 8067 12291
rect 8125 12257 8159 12291
rect 8309 12257 8343 12291
rect 8401 12257 8435 12291
rect 8585 12257 8619 12291
rect 8677 12257 8711 12291
rect 8861 12257 8895 12291
rect 8953 12257 8987 12291
rect 9413 12257 9447 12291
rect 9597 12257 9631 12291
rect 9689 12257 9723 12291
rect 9781 12257 9815 12291
rect 11529 12257 11563 12291
rect 11713 12257 11747 12291
rect 11805 12257 11839 12291
rect 11897 12257 11931 12291
rect 13461 12257 13495 12291
rect 13553 12257 13587 12291
rect 13645 12257 13679 12291
rect 13829 12257 13863 12291
rect 15025 12257 15059 12291
rect 15301 12257 15335 12291
rect 15485 12257 15519 12291
rect 15577 12257 15611 12291
rect 15669 12257 15703 12291
rect 16497 12257 16531 12291
rect 16589 12257 16623 12291
rect 16773 12257 16807 12291
rect 16865 12257 16899 12291
rect 17049 12257 17083 12291
rect 17141 12257 17175 12291
rect 17325 12257 17359 12291
rect 17417 12257 17451 12291
rect 17601 12257 17635 12291
rect 17693 12257 17727 12291
rect 17877 12257 17911 12291
rect 17969 12257 18003 12291
rect 18153 12257 18187 12291
rect 18245 12257 18279 12291
rect 18429 12257 18463 12291
rect 18521 12257 18555 12291
rect 18705 12257 18739 12291
rect 18797 12257 18831 12291
rect 18981 12257 19015 12291
rect 19073 12257 19107 12291
rect 19257 12257 19291 12291
rect 19349 12257 19383 12291
rect 19533 12257 19567 12291
rect 20269 12257 20303 12291
rect 20545 12257 20579 12291
rect 20637 12257 20671 12291
rect 22017 12257 22051 12291
rect 22293 12257 22327 12291
rect 22385 12257 22419 12291
rect 22477 12257 22511 12291
rect 22661 12257 22695 12291
rect 24409 12257 24443 12291
rect 24593 12257 24627 12291
rect 24685 12257 24719 12291
rect 24869 12257 24903 12291
rect 24961 12257 24995 12291
rect 25053 12257 25087 12291
rect 26617 12257 26651 12291
rect 26709 12257 26743 12291
rect 26801 12257 26835 12291
rect 26985 12257 27019 12291
rect 28365 12257 28399 12291
rect 28549 12257 28583 12291
rect 28641 12257 28675 12291
rect 28733 12257 28767 12291
rect 30113 12257 30147 12291
rect 30389 12257 30423 12291
rect 30481 12257 30515 12291
rect 30757 12257 30791 12291
rect 2881 12189 2915 12223
rect 9873 12189 9907 12223
rect 13369 12189 13403 12223
rect 15761 12189 15795 12223
rect 20729 12189 20763 12223
rect 22753 12189 22787 12223
rect 25145 12189 25179 12223
rect 26525 12189 26559 12223
rect 28825 12189 28859 12223
rect 30297 12189 30331 12223
rect 30021 12121 30055 12155
rect 3157 12053 3191 12087
rect 6101 12053 6135 12087
rect 11437 12053 11471 12087
rect 15209 12053 15243 12087
rect 20453 12053 20487 12087
rect 24317 12053 24351 12087
rect 28273 12053 28307 12087
rect 6285 11849 6319 11883
rect 9689 11849 9723 11883
rect 13645 11849 13679 11883
rect 16313 11849 16347 11883
rect 22293 11849 22327 11883
rect 27077 11849 27111 11883
rect 30389 11849 30423 11883
rect 10517 11713 10551 11747
rect 13001 11713 13035 11747
rect 14197 11713 14231 11747
rect 21097 11713 21131 11747
rect 25053 11713 25087 11747
rect 25973 11713 26007 11747
rect 28181 11713 28215 11747
rect 30113 11713 30147 11747
rect 3249 11645 3283 11679
rect 3341 11645 3375 11679
rect 3525 11645 3559 11679
rect 3617 11645 3651 11679
rect 3801 11645 3835 11679
rect 3893 11645 3927 11679
rect 4077 11645 4111 11679
rect 6193 11645 6227 11679
rect 9505 11645 9539 11679
rect 9781 11645 9815 11679
rect 9965 11645 9999 11679
rect 10057 11645 10091 11679
rect 10241 11645 10275 11679
rect 10333 11645 10367 11679
rect 10425 11645 10459 11679
rect 11345 11645 11379 11679
rect 11437 11645 11471 11679
rect 11529 11645 11563 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 13093 11645 13127 11679
rect 13185 11645 13219 11679
rect 13737 11645 13771 11679
rect 13921 11645 13955 11679
rect 14013 11645 14047 11679
rect 14105 11645 14139 11679
rect 15117 11645 15151 11679
rect 15209 11645 15243 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 15669 11645 15703 11679
rect 15761 11645 15795 11679
rect 15945 11645 15979 11679
rect 16037 11645 16071 11679
rect 16221 11645 16255 11679
rect 20361 11645 20395 11679
rect 20453 11645 20487 11679
rect 20545 11645 20579 11679
rect 20729 11645 20763 11679
rect 20821 11645 20855 11679
rect 21005 11645 21039 11679
rect 22385 11645 22419 11679
rect 22569 11645 22603 11679
rect 22661 11645 22695 11679
rect 22845 11645 22879 11679
rect 22937 11645 22971 11679
rect 23121 11645 23155 11679
rect 23213 11645 23247 11679
rect 23397 11645 23431 11679
rect 23489 11645 23523 11679
rect 23949 11645 23983 11679
rect 24041 11645 24075 11679
rect 24225 11645 24259 11679
rect 24317 11645 24351 11679
rect 24501 11645 24535 11679
rect 24593 11645 24627 11679
rect 24777 11645 24811 11679
rect 24869 11645 24903 11679
rect 24961 11645 24995 11679
rect 25789 11645 25823 11679
rect 25881 11645 25915 11679
rect 26157 11645 26191 11679
rect 26249 11645 26283 11679
rect 26433 11645 26467 11679
rect 26525 11645 26559 11679
rect 26709 11645 26743 11679
rect 26801 11645 26835 11679
rect 26985 11645 27019 11679
rect 27997 11645 28031 11679
rect 28273 11645 28307 11679
rect 28365 11645 28399 11679
rect 28457 11645 28491 11679
rect 28641 11645 28675 11679
rect 30205 11645 30239 11679
rect 30481 11645 30515 11679
rect 30665 11645 30699 11679
rect 30757 11645 30791 11679
rect 30941 11645 30975 11679
rect 31033 11645 31067 11679
rect 31125 11645 31159 11679
rect 9413 11577 9447 11611
rect 12357 11577 12391 11611
rect 13277 11577 13311 11611
rect 25697 11577 25731 11611
rect 28733 11577 28767 11611
rect 31217 11577 31251 11611
rect 4169 11509 4203 11543
rect 11253 11509 11287 11543
rect 20269 11509 20303 11543
rect 27905 11509 27939 11543
rect 7573 11305 7607 11339
rect 9689 11305 9723 11339
rect 13277 11305 13311 11339
rect 25513 11305 25547 11339
rect 30665 11305 30699 11339
rect 3433 11237 3467 11271
rect 5273 11237 5307 11271
rect 5917 11237 5951 11271
rect 7849 11237 7883 11271
rect 10241 11237 10275 11271
rect 13829 11237 13863 11271
rect 16221 11237 16255 11271
rect 17693 11237 17727 11271
rect 20729 11237 20763 11271
rect 26065 11237 26099 11271
rect 28273 11237 28307 11271
rect 29285 11237 29319 11271
rect 3525 11169 3559 11203
rect 3617 11169 3651 11203
rect 3709 11169 3743 11203
rect 3893 11169 3927 11203
rect 5365 11169 5399 11203
rect 5457 11169 5491 11203
rect 6009 11169 6043 11203
rect 6101 11169 6135 11203
rect 6193 11169 6227 11203
rect 6377 11169 6411 11203
rect 6469 11169 6503 11203
rect 6653 11169 6687 11203
rect 6745 11169 6779 11203
rect 6929 11169 6963 11203
rect 7021 11169 7055 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 7481 11169 7515 11203
rect 7941 11169 7975 11203
rect 8033 11169 8067 11203
rect 8309 11169 8343 11203
rect 9781 11169 9815 11203
rect 9965 11169 9999 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 11529 11169 11563 11203
rect 11621 11169 11655 11203
rect 11805 11169 11839 11203
rect 13369 11169 13403 11203
rect 13553 11169 13587 11203
rect 13645 11169 13679 11203
rect 13737 11169 13771 11203
rect 14657 11169 14691 11203
rect 14841 11169 14875 11203
rect 14933 11169 14967 11203
rect 15117 11169 15151 11203
rect 15209 11169 15243 11203
rect 15393 11169 15427 11203
rect 15485 11169 15519 11203
rect 15853 11169 15887 11203
rect 16129 11169 16163 11203
rect 17785 11169 17819 11203
rect 17877 11169 17911 11203
rect 18337 11169 18371 11203
rect 18521 11169 18555 11203
rect 18613 11169 18647 11203
rect 18797 11169 18831 11203
rect 18889 11169 18923 11203
rect 19073 11169 19107 11203
rect 19165 11169 19199 11203
rect 19349 11169 19383 11203
rect 19441 11169 19475 11203
rect 19625 11169 19659 11203
rect 19717 11169 19751 11203
rect 19901 11169 19935 11203
rect 19993 11169 20027 11203
rect 20177 11169 20211 11203
rect 20269 11169 20303 11203
rect 20453 11169 20487 11203
rect 20545 11169 20579 11203
rect 20637 11169 20671 11203
rect 20913 11169 20947 11203
rect 22937 11169 22971 11203
rect 25145 11169 25179 11203
rect 25605 11169 25639 11203
rect 25789 11169 25823 11203
rect 25881 11169 25915 11203
rect 25973 11169 26007 11203
rect 27537 11169 27571 11203
rect 27721 11169 27755 11203
rect 27813 11169 27847 11203
rect 27997 11169 28031 11203
rect 28089 11169 28123 11203
rect 28181 11169 28215 11203
rect 29377 11169 29411 11203
rect 29469 11169 29503 11203
rect 29561 11169 29595 11203
rect 29745 11169 29779 11203
rect 29837 11169 29871 11203
rect 30021 11169 30055 11203
rect 30113 11169 30147 11203
rect 30297 11169 30331 11203
rect 30389 11169 30423 11203
rect 30573 11169 30607 11203
rect 8401 11101 8435 11135
rect 15761 11101 15795 11135
rect 18245 11101 18279 11135
rect 23029 11033 23063 11067
rect 3985 10965 4019 10999
rect 5549 10965 5583 10999
rect 8125 10965 8159 10999
rect 11897 10965 11931 10999
rect 14565 10965 14599 10999
rect 17969 10965 18003 10999
rect 21005 10965 21039 10999
rect 25237 10965 25271 10999
rect 27445 10965 27479 10999
rect 5641 10761 5675 10795
rect 6101 10761 6135 10795
rect 9505 10761 9539 10795
rect 13001 10761 13035 10795
rect 16589 10761 16623 10795
rect 20085 10761 20119 10795
rect 25881 10761 25915 10795
rect 29377 10761 29411 10795
rect 4261 10693 4295 10727
rect 28733 10693 28767 10727
rect 3709 10625 3743 10659
rect 5089 10625 5123 10659
rect 8493 10625 8527 10659
rect 11713 10625 11747 10659
rect 16037 10625 16071 10659
rect 17601 10625 17635 10659
rect 21005 10625 21039 10659
rect 26157 10625 26191 10659
rect 27261 10625 27295 10659
rect 29101 10625 29135 10659
rect 3065 10557 3099 10591
rect 3433 10557 3467 10591
rect 3525 10557 3559 10591
rect 3801 10557 3835 10591
rect 3893 10557 3927 10591
rect 3985 10557 4019 10591
rect 4169 10557 4203 10591
rect 5181 10557 5215 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 5549 10557 5583 10591
rect 6009 10557 6043 10591
rect 7757 10557 7791 10591
rect 8033 10557 8067 10591
rect 8401 10557 8435 10591
rect 9597 10557 9631 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 10149 10557 10183 10591
rect 10333 10557 10367 10591
rect 10425 10557 10459 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 10885 10557 10919 10591
rect 10977 10557 11011 10591
rect 11161 10557 11195 10591
rect 11253 10557 11287 10591
rect 11437 10557 11471 10591
rect 11529 10557 11563 10591
rect 11805 10557 11839 10591
rect 11897 10557 11931 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 13369 10557 13403 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 14565 10557 14599 10591
rect 14657 10557 14691 10591
rect 16129 10557 16163 10591
rect 16313 10557 16347 10591
rect 16405 10557 16439 10591
rect 16497 10557 16531 10591
rect 16773 10557 16807 10591
rect 17693 10557 17727 10591
rect 17785 10557 17819 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 20177 10557 20211 10591
rect 21097 10557 21131 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 21465 10557 21499 10591
rect 21557 10557 21591 10591
rect 21741 10557 21775 10591
rect 21833 10557 21867 10591
rect 22017 10557 22051 10591
rect 22109 10557 22143 10591
rect 22293 10557 22327 10591
rect 22385 10557 22419 10591
rect 22569 10557 22603 10591
rect 22661 10557 22695 10591
rect 22845 10557 22879 10591
rect 22937 10557 22971 10591
rect 23121 10557 23155 10591
rect 23213 10557 23247 10591
rect 23397 10557 23431 10591
rect 23857 10557 23891 10591
rect 23949 10557 23983 10591
rect 24133 10557 24167 10591
rect 24409 10557 24443 10591
rect 24501 10557 24535 10591
rect 24685 10557 24719 10591
rect 24961 10557 24995 10591
rect 25053 10557 25087 10591
rect 25237 10557 25271 10591
rect 25329 10557 25363 10591
rect 25513 10557 25547 10591
rect 25973 10557 26007 10591
rect 26065 10557 26099 10591
rect 26801 10557 26835 10591
rect 26985 10557 27019 10591
rect 27077 10557 27111 10591
rect 27353 10557 27387 10591
rect 27445 10557 27479 10591
rect 28825 10557 28859 10591
rect 29193 10557 29227 10591
rect 29285 10557 29319 10591
rect 29561 10557 29595 10591
rect 7941 10489 7975 10523
rect 12265 10489 12299 10523
rect 16865 10489 16899 10523
rect 27537 10489 27571 10523
rect 29653 10489 29687 10523
rect 2973 10421 3007 10455
rect 7665 10421 7699 10455
rect 9781 10421 9815 10455
rect 18153 10421 18187 10455
rect 23489 10421 23523 10455
rect 24225 10421 24259 10455
rect 24777 10421 24811 10455
rect 25605 10421 25639 10455
rect 26709 10421 26743 10455
rect 5365 10217 5399 10251
rect 7481 10217 7515 10251
rect 9873 10217 9907 10251
rect 16405 10217 16439 10251
rect 21649 10217 21683 10251
rect 22845 10217 22879 10251
rect 23581 10217 23615 10251
rect 24409 10217 24443 10251
rect 25145 10217 25179 10251
rect 28825 10217 28859 10251
rect 3893 10149 3927 10183
rect 5917 10149 5951 10183
rect 7757 10149 7791 10183
rect 16957 10149 16991 10183
rect 27353 10149 27387 10183
rect 29653 10149 29687 10183
rect 3157 10081 3191 10115
rect 3249 10081 3283 10115
rect 3341 10081 3375 10115
rect 3525 10081 3559 10115
rect 3617 10081 3651 10115
rect 3801 10081 3835 10115
rect 4905 10081 4939 10115
rect 5181 10081 5215 10115
rect 5457 10081 5491 10115
rect 5825 10081 5859 10115
rect 6101 10081 6135 10115
rect 7573 10081 7607 10115
rect 7665 10081 7699 10115
rect 8125 10081 8159 10115
rect 8217 10081 8251 10115
rect 8493 10081 8527 10115
rect 9781 10081 9815 10115
rect 16497 10081 16531 10115
rect 16681 10081 16715 10115
rect 16773 10081 16807 10115
rect 16865 10081 16899 10115
rect 17877 10081 17911 10115
rect 17969 10081 18003 10115
rect 18061 10081 18095 10115
rect 18245 10081 18279 10115
rect 18337 10081 18371 10115
rect 18521 10081 18555 10115
rect 19809 10081 19843 10115
rect 19901 10081 19935 10115
rect 19993 10081 20027 10115
rect 20177 10081 20211 10115
rect 20269 10081 20303 10115
rect 20453 10081 20487 10115
rect 20545 10081 20579 10115
rect 20729 10081 20763 10115
rect 20821 10081 20855 10115
rect 21281 10081 21315 10115
rect 21373 10081 21407 10115
rect 21557 10081 21591 10115
rect 22937 10081 22971 10115
rect 23673 10081 23707 10115
rect 24225 10081 24259 10115
rect 24317 10081 24351 10115
rect 25237 10081 25271 10115
rect 26617 10081 26651 10115
rect 26709 10081 26743 10115
rect 26801 10081 26835 10115
rect 26985 10081 27019 10115
rect 27077 10081 27111 10115
rect 27261 10081 27295 10115
rect 28917 10081 28951 10115
rect 29101 10081 29135 10115
rect 29193 10081 29227 10115
rect 29377 10081 29411 10115
rect 29469 10081 29503 10115
rect 29561 10081 29595 10115
rect 5089 10013 5123 10047
rect 8585 10013 8619 10047
rect 17785 10013 17819 10047
rect 19717 10013 19751 10047
rect 24133 10013 24167 10047
rect 6193 9945 6227 9979
rect 8309 9945 8343 9979
rect 3065 9877 3099 9911
rect 4813 9877 4847 9911
rect 8033 9877 8067 9911
rect 18613 9877 18647 9911
rect 26525 9877 26559 9911
rect 5181 9673 5215 9707
rect 16681 9673 16715 9707
rect 20177 9673 20211 9707
rect 29101 9673 29135 9707
rect 15117 9605 15151 9639
rect 4905 9537 4939 9571
rect 10977 9537 11011 9571
rect 14841 9537 14875 9571
rect 18337 9537 18371 9571
rect 28733 9537 28767 9571
rect 3249 9469 3283 9503
rect 3341 9469 3375 9503
rect 3525 9469 3559 9503
rect 3617 9469 3651 9503
rect 3801 9469 3835 9503
rect 3893 9469 3927 9503
rect 4077 9469 4111 9503
rect 4537 9469 4571 9503
rect 4813 9469 4847 9503
rect 5273 9469 5307 9503
rect 5365 9469 5399 9503
rect 7941 9469 7975 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 8677 9469 8711 9503
rect 8769 9469 8803 9503
rect 8953 9469 8987 9503
rect 9045 9469 9079 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 9505 9469 9539 9503
rect 9597 9469 9631 9503
rect 9781 9469 9815 9503
rect 9873 9469 9907 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 10333 9469 10367 9503
rect 10425 9469 10459 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 10885 9469 10919 9503
rect 11437 9469 11471 9503
rect 11529 9469 11563 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 13001 9469 13035 9503
rect 13185 9469 13219 9503
rect 13277 9469 13311 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 13921 9469 13955 9503
rect 14013 9469 14047 9503
rect 14197 9469 14231 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 14749 9469 14783 9503
rect 15209 9469 15243 9503
rect 15301 9469 15335 9503
rect 15577 9469 15611 9503
rect 16773 9469 16807 9503
rect 16957 9469 16991 9503
rect 17049 9469 17083 9503
rect 17233 9469 17267 9503
rect 17325 9469 17359 9503
rect 17417 9469 17451 9503
rect 18429 9469 18463 9503
rect 18705 9469 18739 9503
rect 18797 9469 18831 9503
rect 18981 9469 19015 9503
rect 19073 9469 19107 9503
rect 19257 9469 19291 9503
rect 19349 9469 19383 9503
rect 19533 9469 19567 9503
rect 19625 9469 19659 9503
rect 19809 9469 19843 9503
rect 19901 9469 19935 9503
rect 20085 9469 20119 9503
rect 22293 9469 22327 9503
rect 22477 9469 22511 9503
rect 22569 9469 22603 9503
rect 22753 9469 22787 9503
rect 22845 9469 22879 9503
rect 23029 9469 23063 9503
rect 23121 9469 23155 9503
rect 23213 9469 23247 9503
rect 26525 9469 26559 9503
rect 26617 9469 26651 9503
rect 26709 9469 26743 9503
rect 26893 9469 26927 9503
rect 26985 9469 27019 9503
rect 27169 9469 27203 9503
rect 28825 9469 28859 9503
rect 29193 9469 29227 9503
rect 29377 9469 29411 9503
rect 29469 9469 29503 9503
rect 29561 9469 29595 9503
rect 4629 9401 4663 9435
rect 5457 9401 5491 9435
rect 7849 9401 7883 9435
rect 8493 9401 8527 9435
rect 11621 9401 11655 9435
rect 12725 9401 12759 9435
rect 15393 9401 15427 9435
rect 17509 9401 17543 9435
rect 23305 9401 23339 9435
rect 27261 9401 27295 9435
rect 29653 9401 29687 9435
rect 4169 9333 4203 9367
rect 8125 9333 8159 9367
rect 11345 9333 11379 9367
rect 15669 9333 15703 9367
rect 22201 9333 22235 9367
rect 26433 9333 26467 9367
rect 4537 9129 4571 9163
rect 8677 9129 8711 9163
rect 13001 9129 13035 9163
rect 17141 9129 17175 9163
rect 23213 9129 23247 9163
rect 28825 9129 28859 9163
rect 4813 9061 4847 9095
rect 12633 9061 12667 9095
rect 15209 9061 15243 9095
rect 29653 9061 29687 9095
rect 3617 8993 3651 9027
rect 3709 8993 3743 9027
rect 4353 8993 4387 9027
rect 4445 8993 4479 9027
rect 4721 8993 4755 9027
rect 7481 8993 7515 9027
rect 8585 8993 8619 9027
rect 11345 8993 11379 9027
rect 11437 8993 11471 9027
rect 11529 8993 11563 9027
rect 11713 8993 11747 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 12081 8993 12115 9027
rect 12265 8993 12299 9027
rect 12357 8993 12391 9027
rect 12541 8993 12575 9027
rect 13093 8993 13127 9027
rect 13185 8993 13219 9027
rect 15025 8993 15059 9027
rect 15301 8993 15335 9027
rect 15393 8993 15427 9027
rect 15485 8993 15519 9027
rect 15669 8993 15703 9027
rect 17233 8993 17267 9027
rect 17417 8993 17451 9027
rect 17509 8993 17543 9027
rect 17693 8993 17727 9027
rect 17785 8993 17819 9027
rect 17877 8993 17911 9027
rect 19073 8993 19107 9027
rect 19533 8993 19567 9027
rect 19717 8993 19751 9027
rect 19809 8993 19843 9027
rect 19993 8993 20027 9027
rect 20085 8993 20119 9027
rect 20269 8993 20303 9027
rect 20361 8993 20395 9027
rect 20545 8993 20579 9027
rect 20637 8993 20671 9027
rect 20821 8993 20855 9027
rect 20913 8993 20947 9027
rect 21373 8993 21407 9027
rect 21465 8993 21499 9027
rect 21649 8993 21683 9027
rect 21741 8993 21775 9027
rect 21925 8993 21959 9027
rect 22017 8993 22051 9027
rect 22201 8993 22235 9027
rect 22293 8993 22327 9027
rect 22385 8993 22419 9027
rect 22661 8993 22695 9027
rect 23305 8993 23339 9027
rect 23489 8993 23523 9027
rect 23581 8993 23615 9027
rect 23765 8993 23799 9027
rect 23857 8993 23891 9027
rect 24041 8993 24075 9027
rect 24133 8993 24167 9027
rect 24317 8993 24351 9027
rect 24409 8993 24443 9027
rect 24501 8993 24535 9027
rect 26525 8993 26559 9027
rect 26617 8993 26651 9027
rect 26801 8993 26835 9027
rect 26893 8993 26927 9027
rect 27077 8993 27111 9027
rect 28917 8993 28951 9027
rect 29101 8993 29135 9027
rect 29193 8993 29227 9027
rect 29377 8993 29411 9027
rect 29469 8993 29503 9027
rect 29561 8993 29595 9027
rect 3525 8925 3559 8959
rect 4261 8925 4295 8959
rect 11253 8925 11287 8959
rect 13277 8925 13311 8959
rect 15761 8925 15795 8959
rect 17969 8925 18003 8959
rect 22477 8925 22511 8959
rect 24593 8925 24627 8959
rect 3801 8857 3835 8891
rect 7573 8789 7607 8823
rect 14933 8789 14967 8823
rect 18981 8789 19015 8823
rect 19441 8789 19475 8823
rect 22753 8789 22787 8823
rect 27169 8789 27203 8823
rect 11529 8585 11563 8619
rect 17233 8585 17267 8619
rect 18981 8585 19015 8619
rect 21833 8585 21867 8619
rect 24041 8585 24075 8619
rect 29377 8585 29411 8619
rect 19809 8517 19843 8551
rect 16957 8449 16991 8483
rect 7389 8381 7423 8415
rect 7665 8381 7699 8415
rect 7849 8381 7883 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 8217 8381 8251 8415
rect 8677 8381 8711 8415
rect 8953 8381 8987 8415
rect 9137 8381 9171 8415
rect 9229 8381 9263 8415
rect 9413 8381 9447 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 9781 8381 9815 8415
rect 9965 8381 9999 8415
rect 10057 8381 10091 8415
rect 10241 8381 10275 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 10609 8381 10643 8415
rect 10701 8381 10735 8415
rect 11437 8381 11471 8415
rect 15117 8381 15151 8415
rect 15209 8381 15243 8415
rect 15393 8381 15427 8415
rect 15485 8381 15519 8415
rect 15669 8381 15703 8415
rect 15761 8381 15795 8415
rect 15945 8381 15979 8415
rect 17049 8381 17083 8415
rect 17325 8381 17359 8415
rect 17509 8381 17543 8415
rect 17601 8381 17635 8415
rect 17693 8381 17727 8415
rect 19073 8381 19107 8415
rect 19349 8381 19383 8415
rect 19441 8381 19475 8415
rect 19533 8381 19567 8415
rect 19717 8381 19751 8415
rect 21925 8381 21959 8415
rect 24133 8381 24167 8415
rect 24317 8381 24351 8415
rect 24409 8381 24443 8415
rect 24501 8381 24535 8415
rect 26709 8381 26743 8415
rect 26801 8381 26835 8415
rect 26893 8381 26927 8415
rect 27077 8381 27111 8415
rect 27169 8381 27203 8415
rect 27353 8381 27387 8415
rect 27445 8381 27479 8415
rect 27629 8381 27663 8415
rect 27721 8381 27755 8415
rect 27905 8381 27939 8415
rect 27997 8381 28031 8415
rect 28181 8381 28215 8415
rect 28273 8381 28307 8415
rect 28457 8381 28491 8415
rect 28549 8381 28583 8415
rect 29009 8381 29043 8415
rect 29285 8381 29319 8415
rect 10793 8313 10827 8347
rect 17785 8313 17819 8347
rect 19257 8313 19291 8347
rect 24593 8313 24627 8347
rect 26617 8313 26651 8347
rect 7297 8245 7331 8279
rect 7573 8245 7607 8279
rect 8585 8245 8619 8279
rect 8861 8245 8895 8279
rect 16037 8245 16071 8279
rect 29101 8245 29135 8279
rect 7573 8041 7607 8075
rect 9137 8041 9171 8075
rect 10701 8041 10735 8075
rect 17233 8041 17267 8075
rect 24133 8041 24167 8075
rect 28733 8041 28767 8075
rect 7849 7973 7883 8007
rect 13737 7973 13771 8007
rect 16221 7973 16255 8007
rect 7481 7905 7515 7939
rect 7757 7905 7791 7939
rect 8033 7905 8067 7939
rect 8125 7905 8159 7939
rect 8309 7905 8343 7939
rect 8585 7905 8619 7939
rect 9045 7905 9079 7939
rect 10793 7905 10827 7939
rect 11345 7905 11379 7939
rect 11529 7905 11563 7939
rect 11621 7905 11655 7939
rect 11805 7905 11839 7939
rect 11897 7905 11931 7939
rect 12081 7905 12115 7939
rect 12173 7905 12207 7939
rect 12357 7905 12391 7939
rect 12449 7905 12483 7939
rect 12633 7905 12667 7939
rect 12725 7905 12759 7939
rect 12909 7905 12943 7939
rect 13001 7905 13035 7939
rect 13185 7905 13219 7939
rect 13277 7905 13311 7939
rect 13553 7905 13587 7939
rect 13645 7905 13679 7939
rect 15117 7905 15151 7939
rect 15393 7905 15427 7939
rect 15485 7905 15519 7939
rect 15577 7905 15611 7939
rect 15761 7905 15795 7939
rect 15853 7905 15887 7939
rect 16129 7905 16163 7939
rect 17325 7905 17359 7939
rect 17509 7905 17543 7939
rect 17601 7905 17635 7939
rect 17785 7905 17819 7939
rect 17877 7905 17911 7939
rect 18061 7905 18095 7939
rect 18153 7905 18187 7939
rect 18337 7905 18371 7939
rect 18429 7905 18463 7939
rect 18613 7905 18647 7939
rect 18705 7905 18739 7939
rect 18889 7905 18923 7939
rect 18981 7905 19015 7939
rect 20361 7905 20395 7939
rect 20453 7905 20487 7939
rect 20545 7905 20579 7939
rect 20729 7905 20763 7939
rect 20821 7905 20855 7939
rect 21281 7905 21315 7939
rect 21373 7905 21407 7939
rect 21557 7905 21591 7939
rect 21649 7905 21683 7939
rect 21833 7905 21867 7939
rect 21925 7905 21959 7939
rect 22109 7905 22143 7939
rect 22201 7905 22235 7939
rect 22385 7905 22419 7939
rect 22661 7905 22695 7939
rect 22753 7905 22787 7939
rect 22937 7905 22971 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 23489 7905 23523 7939
rect 24225 7905 24259 7939
rect 24409 7905 24443 7939
rect 24501 7905 24535 7939
rect 24685 7905 24719 7939
rect 24777 7905 24811 7939
rect 24961 7905 24995 7939
rect 25053 7905 25087 7939
rect 25237 7905 25271 7939
rect 25329 7905 25363 7939
rect 25513 7905 25547 7939
rect 25605 7905 25639 7939
rect 25789 7905 25823 7939
rect 25881 7905 25915 7939
rect 25973 7905 26007 7939
rect 28825 7905 28859 7939
rect 29009 7905 29043 7939
rect 29101 7905 29135 7939
rect 8677 7837 8711 7871
rect 13461 7837 13495 7871
rect 15301 7837 15335 7871
rect 20269 7837 20303 7871
rect 26065 7837 26099 7871
rect 23581 7769 23615 7803
rect 8401 7701 8435 7735
rect 11253 7701 11287 7735
rect 15025 7701 15059 7735
rect 22477 7701 22511 7735
rect 23305 7701 23339 7735
rect 11253 7497 11287 7531
rect 13645 7497 13679 7531
rect 20545 7497 20579 7531
rect 21833 7497 21867 7531
rect 25329 7497 25363 7531
rect 17233 7429 17267 7463
rect 19993 7429 20027 7463
rect 7573 7361 7607 7395
rect 9597 7361 9631 7395
rect 11529 7361 11563 7395
rect 14197 7361 14231 7395
rect 20269 7361 20303 7395
rect 22661 7361 22695 7395
rect 22937 7361 22971 7395
rect 25881 7361 25915 7395
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 7389 7293 7423 7327
rect 7665 7293 7699 7327
rect 7757 7293 7791 7327
rect 7849 7293 7883 7327
rect 8033 7293 8067 7327
rect 8125 7293 8159 7327
rect 8401 7293 8435 7327
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 8953 7293 8987 7327
rect 9045 7293 9079 7327
rect 9229 7293 9263 7327
rect 9321 7293 9355 7327
rect 9505 7293 9539 7327
rect 9965 7293 9999 7327
rect 10057 7293 10091 7327
rect 11345 7293 11379 7327
rect 11437 7293 11471 7327
rect 13737 7293 13771 7327
rect 13921 7293 13955 7327
rect 14013 7293 14047 7327
rect 14105 7293 14139 7327
rect 15209 7293 15243 7327
rect 15301 7293 15335 7327
rect 15485 7293 15519 7327
rect 15577 7293 15611 7327
rect 15761 7293 15795 7327
rect 17141 7293 17175 7327
rect 17417 7293 17451 7327
rect 17509 7293 17543 7327
rect 17693 7293 17727 7327
rect 18061 7293 18095 7327
rect 19809 7293 19843 7327
rect 20085 7293 20119 7327
rect 20177 7293 20211 7327
rect 20453 7293 20487 7327
rect 21925 7293 21959 7327
rect 22753 7293 22787 7327
rect 23029 7293 23063 7327
rect 23121 7293 23155 7327
rect 23213 7293 23247 7327
rect 23397 7293 23431 7327
rect 25421 7293 25455 7327
rect 25605 7293 25639 7327
rect 25697 7293 25731 7327
rect 25789 7293 25823 7327
rect 10149 7225 10183 7259
rect 19717 7225 19751 7259
rect 7021 7157 7055 7191
rect 9873 7157 9907 7191
rect 15853 7157 15887 7191
rect 17785 7157 17819 7191
rect 18153 7157 18187 7191
rect 23489 7157 23523 7191
rect 7849 6953 7883 6987
rect 17141 6953 17175 6987
rect 19809 6953 19843 6987
rect 25329 6953 25363 6987
rect 6653 6817 6687 6851
rect 6837 6817 6871 6851
rect 6929 6817 6963 6851
rect 7113 6817 7147 6851
rect 7205 6817 7239 6851
rect 7757 6817 7791 6851
rect 9873 6817 9907 6851
rect 9965 6817 9999 6851
rect 10057 6817 10091 6851
rect 10241 6817 10275 6851
rect 10333 6817 10367 6851
rect 10517 6817 10551 6851
rect 13461 6817 13495 6851
rect 13737 6817 13771 6851
rect 13921 6817 13955 6851
rect 14013 6817 14047 6851
rect 14197 6817 14231 6851
rect 14289 6817 14323 6851
rect 14473 6817 14507 6851
rect 14565 6817 14599 6851
rect 14749 6817 14783 6851
rect 14841 6817 14875 6851
rect 15209 6817 15243 6851
rect 15301 6817 15335 6851
rect 15945 6817 15979 6851
rect 16221 6817 16255 6851
rect 16313 6817 16347 6851
rect 16497 6817 16531 6851
rect 16589 6817 16623 6851
rect 16957 6817 16991 6851
rect 17049 6817 17083 6851
rect 17325 6817 17359 6851
rect 17785 6817 17819 6851
rect 17877 6817 17911 6851
rect 18245 6817 18279 6851
rect 18337 6817 18371 6851
rect 18613 6817 18647 6851
rect 18705 6817 18739 6851
rect 18889 6817 18923 6851
rect 18981 6817 19015 6851
rect 19165 6817 19199 6851
rect 19257 6817 19291 6851
rect 19441 6817 19475 6851
rect 19533 6817 19567 6851
rect 19901 6817 19935 6851
rect 19993 6817 20027 6851
rect 22017 6817 22051 6851
rect 22201 6817 22235 6851
rect 22293 6817 22327 6851
rect 22477 6817 22511 6851
rect 22569 6817 22603 6851
rect 22753 6817 22787 6851
rect 22845 6817 22879 6851
rect 23121 6817 23155 6851
rect 23213 6817 23247 6851
rect 25421 6817 25455 6851
rect 25605 6817 25639 6851
rect 25697 6817 25731 6851
rect 25881 6817 25915 6851
rect 25973 6817 26007 6851
rect 26065 6817 26099 6851
rect 10609 6749 10643 6783
rect 13369 6749 13403 6783
rect 15117 6749 15151 6783
rect 15853 6749 15887 6783
rect 16865 6749 16899 6783
rect 20085 6749 20119 6783
rect 23029 6749 23063 6783
rect 26157 6749 26191 6783
rect 15393 6681 15427 6715
rect 17417 6681 17451 6715
rect 23305 6681 23339 6715
rect 6561 6613 6595 6647
rect 9781 6613 9815 6647
rect 13645 6613 13679 6647
rect 21925 6613 21959 6647
rect 7205 6409 7239 6443
rect 13737 6409 13771 6443
rect 16221 6409 16255 6443
rect 25329 6409 25363 6443
rect 21557 6341 21591 6375
rect 6653 6273 6687 6307
rect 8493 6273 8527 6307
rect 11621 6273 11655 6307
rect 13093 6273 13127 6307
rect 16497 6273 16531 6307
rect 22385 6273 22419 6307
rect 5917 6205 5951 6239
rect 6193 6205 6227 6239
rect 6377 6205 6411 6239
rect 6469 6205 6503 6239
rect 6561 6205 6595 6239
rect 7297 6205 7331 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 7849 6205 7883 6239
rect 8033 6205 8067 6239
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 10057 6205 10091 6239
rect 10149 6205 10183 6239
rect 10333 6205 10367 6239
rect 11161 6205 11195 6239
rect 11253 6205 11287 6239
rect 11713 6205 11747 6239
rect 11805 6205 11839 6239
rect 11897 6205 11931 6239
rect 12081 6205 12115 6239
rect 12173 6205 12207 6239
rect 12357 6205 12391 6239
rect 12909 6205 12943 6239
rect 13001 6205 13035 6239
rect 13645 6205 13679 6239
rect 16037 6205 16071 6239
rect 16313 6205 16347 6239
rect 16405 6205 16439 6239
rect 16681 6205 16715 6239
rect 21649 6205 21683 6239
rect 21925 6205 21959 6239
rect 22017 6205 22051 6239
rect 22109 6205 22143 6239
rect 22293 6205 22327 6239
rect 22569 6205 22603 6239
rect 25421 6205 25455 6239
rect 25605 6205 25639 6239
rect 25697 6205 25731 6239
rect 25881 6205 25915 6239
rect 25973 6205 26007 6239
rect 26065 6205 26099 6239
rect 6101 6137 6135 6171
rect 11069 6137 11103 6171
rect 12449 6137 12483 6171
rect 15945 6137 15979 6171
rect 21833 6137 21867 6171
rect 26157 6137 26191 6171
rect 5825 6069 5859 6103
rect 10425 6069 10459 6103
rect 11345 6069 11379 6103
rect 12817 6069 12851 6103
rect 16773 6069 16807 6103
rect 22661 6069 22695 6103
rect 8217 5865 8251 5899
rect 11345 5865 11379 5899
rect 11897 5865 11931 5899
rect 15853 5865 15887 5899
rect 25329 5865 25363 5899
rect 6653 5797 6687 5831
rect 9597 5797 9631 5831
rect 11621 5797 11655 5831
rect 12541 5797 12575 5831
rect 13921 5797 13955 5831
rect 16497 5797 16531 5831
rect 25881 5797 25915 5831
rect 5641 5729 5675 5763
rect 5825 5729 5859 5763
rect 6469 5729 6503 5763
rect 6561 5729 6595 5763
rect 8309 5729 8343 5763
rect 8493 5729 8527 5763
rect 8585 5729 8619 5763
rect 8861 5729 8895 5763
rect 9045 5729 9079 5763
rect 9137 5729 9171 5763
rect 9229 5729 9263 5763
rect 9505 5729 9539 5763
rect 9965 5729 9999 5763
rect 10149 5729 10183 5763
rect 10241 5729 10275 5763
rect 10333 5729 10367 5763
rect 10425 5729 10459 5763
rect 10609 5729 10643 5763
rect 11161 5729 11195 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 11805 5729 11839 5763
rect 12633 5729 12667 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 13001 5729 13035 5763
rect 13093 5729 13127 5763
rect 13277 5729 13311 5763
rect 13369 5729 13403 5763
rect 13553 5729 13587 5763
rect 13645 5729 13679 5763
rect 13829 5729 13863 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 15945 5729 15979 5763
rect 16221 5729 16255 5763
rect 16313 5729 16347 5763
rect 16405 5729 16439 5763
rect 17325 5729 17359 5763
rect 17509 5729 17543 5763
rect 17601 5729 17635 5763
rect 17785 5729 17819 5763
rect 17877 5729 17911 5763
rect 18061 5729 18095 5763
rect 18153 5729 18187 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 18613 5729 18647 5763
rect 18705 5729 18739 5763
rect 18889 5729 18923 5763
rect 18981 5729 19015 5763
rect 19165 5729 19199 5763
rect 19257 5729 19291 5763
rect 19349 5729 19383 5763
rect 19809 5729 19843 5763
rect 19993 5729 20027 5763
rect 20085 5729 20119 5763
rect 20269 5729 20303 5763
rect 20361 5729 20395 5763
rect 20453 5729 20487 5763
rect 20729 5729 20763 5763
rect 22017 5729 22051 5763
rect 22109 5729 22143 5763
rect 22201 5729 22235 5763
rect 22385 5729 22419 5763
rect 22477 5729 22511 5763
rect 22661 5729 22695 5763
rect 24961 5729 24995 5763
rect 25421 5729 25455 5763
rect 25605 5729 25639 5763
rect 25697 5729 25731 5763
rect 25789 5729 25823 5763
rect 5917 5661 5951 5695
rect 8769 5661 8803 5695
rect 9873 5661 9907 5695
rect 11069 5661 11103 5695
rect 14565 5661 14599 5695
rect 19441 5661 19475 5695
rect 20545 5661 20579 5695
rect 21925 5661 21959 5695
rect 25053 5661 25087 5695
rect 5549 5593 5583 5627
rect 9321 5593 9355 5627
rect 10701 5593 10735 5627
rect 6377 5525 6411 5559
rect 14289 5525 14323 5559
rect 17233 5525 17267 5559
rect 19717 5525 19751 5559
rect 20821 5525 20855 5559
rect 22753 5525 22787 5559
rect 9045 5321 9079 5355
rect 15945 5321 15979 5355
rect 18797 5321 18831 5355
rect 20269 5321 20303 5355
rect 6837 5253 6871 5287
rect 14381 5253 14415 5287
rect 19901 5253 19935 5287
rect 7113 5185 7147 5219
rect 21373 5185 21407 5219
rect 22385 5185 22419 5219
rect 6469 5117 6503 5151
rect 6929 5117 6963 5151
rect 7021 5117 7055 5151
rect 7297 5117 7331 5151
rect 9137 5117 9171 5151
rect 9321 5117 9355 5151
rect 9413 5117 9447 5151
rect 9505 5117 9539 5151
rect 14289 5117 14323 5151
rect 14749 5117 14783 5151
rect 14841 5117 14875 5151
rect 15117 5117 15151 5151
rect 16037 5117 16071 5151
rect 16221 5117 16255 5151
rect 16313 5117 16347 5151
rect 16497 5117 16531 5151
rect 16589 5117 16623 5151
rect 16773 5117 16807 5151
rect 16865 5117 16899 5151
rect 17049 5117 17083 5151
rect 17141 5117 17175 5151
rect 18889 5117 18923 5151
rect 19993 5117 20027 5151
rect 20361 5117 20395 5151
rect 20545 5117 20579 5151
rect 20637 5117 20671 5151
rect 20821 5117 20855 5151
rect 20913 5117 20947 5151
rect 21097 5117 21131 5151
rect 21189 5117 21223 5151
rect 21281 5117 21315 5151
rect 22477 5117 22511 5151
rect 22569 5117 22603 5151
rect 22661 5117 22695 5151
rect 22845 5117 22879 5151
rect 22937 5117 22971 5151
rect 23121 5117 23155 5151
rect 23213 5117 23247 5151
rect 23397 5117 23431 5151
rect 23489 5117 23523 5151
rect 23857 5117 23891 5151
rect 23949 5117 23983 5151
rect 24133 5117 24167 5151
rect 24225 5117 24259 5151
rect 24409 5117 24443 5151
rect 24501 5117 24535 5151
rect 24685 5117 24719 5151
rect 24777 5117 24811 5151
rect 24961 5117 24995 5151
rect 25237 5117 25271 5151
rect 25329 5117 25363 5151
rect 25513 5117 25547 5151
rect 6561 5049 6595 5083
rect 9597 5049 9631 5083
rect 14657 5049 14691 5083
rect 15209 5049 15243 5083
rect 7389 4981 7423 5015
rect 14933 4981 14967 5015
rect 25053 4981 25087 5015
rect 25605 4981 25639 5015
rect 8953 4777 8987 4811
rect 21005 4777 21039 4811
rect 24409 4777 24443 4811
rect 24961 4777 24995 4811
rect 8677 4709 8711 4743
rect 13461 4709 13495 4743
rect 15301 4709 15335 4743
rect 7021 4641 7055 4675
rect 7113 4641 7147 4675
rect 7205 4641 7239 4675
rect 7389 4641 7423 4675
rect 7481 4641 7515 4675
rect 7665 4641 7699 4675
rect 8585 4641 8619 4675
rect 9045 4641 9079 4675
rect 9229 4641 9263 4675
rect 9321 4641 9355 4675
rect 9413 4641 9447 4675
rect 11437 4641 11471 4675
rect 11621 4641 11655 4675
rect 11713 4641 11747 4675
rect 11989 4641 12023 4675
rect 12173 4641 12207 4675
rect 12265 4641 12299 4675
rect 12449 4641 12483 4675
rect 12541 4641 12575 4675
rect 12725 4641 12759 4675
rect 12817 4641 12851 4675
rect 13001 4641 13035 4675
rect 13093 4641 13127 4675
rect 13553 4641 13587 4675
rect 13737 4641 13771 4675
rect 13829 4641 13863 4675
rect 13921 4641 13955 4675
rect 14933 4641 14967 4675
rect 15025 4641 15059 4675
rect 15209 4641 15243 4675
rect 15761 4641 15795 4675
rect 16129 4641 16163 4675
rect 17417 4641 17451 4675
rect 17509 4641 17543 4675
rect 17693 4641 17727 4675
rect 17785 4641 17819 4675
rect 17969 4641 18003 4675
rect 18061 4641 18095 4675
rect 18245 4641 18279 4675
rect 18337 4641 18371 4675
rect 18521 4641 18555 4675
rect 18613 4641 18647 4675
rect 18797 4641 18831 4675
rect 18889 4641 18923 4675
rect 19073 4641 19107 4675
rect 19165 4641 19199 4675
rect 19349 4641 19383 4675
rect 19441 4641 19475 4675
rect 19625 4641 19659 4675
rect 19717 4641 19751 4675
rect 19901 4641 19935 4675
rect 21097 4641 21131 4675
rect 21373 4641 21407 4675
rect 21465 4641 21499 4675
rect 21649 4641 21683 4675
rect 21741 4641 21775 4675
rect 21833 4641 21867 4675
rect 24501 4641 24535 4675
rect 25053 4641 25087 4675
rect 6929 4573 6963 4607
rect 9505 4573 9539 4607
rect 14013 4573 14047 4607
rect 16221 4573 16255 4607
rect 21925 4573 21959 4607
rect 7757 4437 7791 4471
rect 11345 4437 11379 4471
rect 11897 4437 11931 4471
rect 15669 4437 15703 4471
rect 19993 4437 20027 4471
rect 8677 4233 8711 4267
rect 12173 4233 12207 4267
rect 17509 4233 17543 4267
rect 21373 4233 21407 4267
rect 7481 4097 7515 4131
rect 8125 4097 8159 4131
rect 6745 4029 6779 4063
rect 7021 4029 7055 4063
rect 7113 4029 7147 4063
rect 7205 4029 7239 4063
rect 7389 4029 7423 4063
rect 8217 4029 8251 4063
rect 8769 4029 8803 4063
rect 8953 4029 8987 4063
rect 9045 4029 9079 4063
rect 9137 4029 9171 4063
rect 10241 4029 10275 4063
rect 10425 4029 10459 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 10977 4029 11011 4063
rect 11069 4029 11103 4063
rect 11253 4029 11287 4063
rect 11345 4029 11379 4063
rect 11437 4029 11471 4063
rect 12081 4029 12115 4063
rect 13921 4029 13955 4063
rect 14105 4029 14139 4063
rect 14197 4029 14231 4063
rect 14381 4029 14415 4063
rect 14473 4029 14507 4063
rect 14657 4029 14691 4063
rect 14749 4029 14783 4063
rect 14933 4029 14967 4063
rect 15025 4029 15059 4063
rect 15209 4029 15243 4063
rect 15301 4029 15335 4063
rect 15485 4029 15519 4063
rect 15577 4029 15611 4063
rect 15669 4029 15703 4063
rect 15761 4029 15795 4063
rect 15945 4029 15979 4063
rect 16037 4029 16071 4063
rect 16221 4029 16255 4063
rect 17601 4029 17635 4063
rect 17785 4029 17819 4063
rect 17877 4029 17911 4063
rect 17969 4029 18003 4063
rect 19625 4029 19659 4063
rect 19717 4029 19751 4063
rect 19809 4029 19843 4063
rect 19993 4029 20027 4063
rect 20085 4029 20119 4063
rect 20269 4029 20303 4063
rect 21465 4029 21499 4063
rect 21649 4029 21683 4063
rect 21741 4029 21775 4063
rect 21925 4029 21959 4063
rect 22017 4029 22051 4063
rect 22201 4029 22235 4063
rect 22293 4029 22327 4063
rect 22477 4029 22511 4063
rect 22569 4029 22603 4063
rect 22753 4029 22787 4063
rect 22845 4029 22879 4063
rect 23029 4029 23063 4063
rect 23121 4029 23155 4063
rect 23305 4029 23339 4063
rect 23397 4029 23431 4063
rect 23581 4029 23615 4063
rect 23673 4029 23707 4063
rect 23949 4029 23983 4063
rect 24041 4029 24075 4063
rect 24225 4029 24259 4063
rect 24317 4029 24351 4063
rect 24501 4029 24535 4063
rect 24593 4029 24627 4063
rect 24777 4029 24811 4063
rect 24869 4029 24903 4063
rect 24961 4029 24995 4063
rect 25237 4029 25271 4063
rect 25697 4029 25731 4063
rect 25789 4029 25823 4063
rect 26249 4029 26283 4063
rect 26433 4029 26467 4063
rect 26525 4029 26559 4063
rect 26709 4029 26743 4063
rect 26801 4029 26835 4063
rect 26893 4029 26927 4063
rect 6929 3961 6963 3995
rect 9229 3961 9263 3995
rect 11529 3961 11563 3995
rect 16313 3961 16347 3995
rect 18061 3961 18095 3995
rect 19533 3961 19567 3995
rect 25053 3961 25087 3995
rect 25881 3961 25915 3995
rect 26985 3961 27019 3995
rect 6653 3893 6687 3927
rect 10149 3893 10183 3927
rect 13829 3893 13863 3927
rect 20361 3893 20395 3927
rect 25329 3893 25363 3927
rect 25605 3893 25639 3927
rect 26157 3893 26191 3927
rect 8309 3689 8343 3723
rect 13921 3689 13955 3723
rect 17325 3689 17359 3723
rect 20453 3689 20487 3723
rect 24409 3689 24443 3723
rect 24685 3689 24719 3723
rect 25237 3689 25271 3723
rect 26525 3689 26559 3723
rect 10609 3621 10643 3655
rect 27629 3621 27663 3655
rect 6745 3553 6779 3587
rect 6837 3553 6871 3587
rect 7021 3553 7055 3587
rect 7113 3553 7147 3587
rect 7297 3553 7331 3587
rect 7389 3553 7423 3587
rect 7573 3553 7607 3587
rect 8401 3553 8435 3587
rect 8677 3553 8711 3587
rect 8861 3553 8895 3587
rect 8953 3553 8987 3587
rect 9137 3553 9171 3587
rect 9229 3553 9263 3587
rect 9413 3553 9447 3587
rect 9505 3553 9539 3587
rect 9689 3553 9723 3587
rect 9781 3553 9815 3587
rect 9965 3553 9999 3587
rect 10057 3553 10091 3587
rect 10241 3553 10275 3587
rect 10333 3553 10367 3587
rect 10517 3553 10551 3587
rect 12725 3553 12759 3587
rect 13277 3553 13311 3587
rect 13829 3553 13863 3587
rect 17417 3553 17451 3587
rect 17601 3553 17635 3587
rect 17693 3553 17727 3587
rect 17877 3553 17911 3587
rect 17969 3553 18003 3587
rect 18061 3553 18095 3587
rect 19441 3553 19475 3587
rect 19625 3553 19659 3587
rect 19717 3553 19751 3587
rect 19993 3553 20027 3587
rect 20085 3553 20119 3587
rect 20177 3553 20211 3587
rect 20361 3553 20395 3587
rect 24501 3553 24535 3587
rect 24777 3553 24811 3587
rect 25329 3553 25363 3587
rect 26617 3553 26651 3587
rect 26801 3553 26835 3587
rect 26893 3553 26927 3587
rect 27077 3553 27111 3587
rect 27169 3553 27203 3587
rect 27353 3553 27387 3587
rect 27445 3553 27479 3587
rect 27537 3553 27571 3587
rect 18153 3485 18187 3519
rect 19901 3485 19935 3519
rect 7665 3349 7699 3383
rect 8585 3349 8619 3383
rect 12817 3349 12851 3383
rect 13369 3349 13403 3383
rect 19349 3349 19383 3383
rect 8769 3145 8803 3179
rect 12633 3145 12667 3179
rect 13001 3145 13035 3179
rect 17693 3145 17727 3179
rect 26709 3145 26743 3179
rect 19257 3077 19291 3111
rect 6561 3009 6595 3043
rect 7113 3009 7147 3043
rect 11529 3009 11563 3043
rect 15761 3009 15795 3043
rect 18981 3009 19015 3043
rect 19809 3009 19843 3043
rect 26433 3009 26467 3043
rect 6653 2941 6687 2975
rect 6837 2941 6871 2975
rect 6929 2941 6963 2975
rect 7021 2941 7055 2975
rect 7573 2941 7607 2975
rect 7665 2941 7699 2975
rect 8677 2941 8711 2975
rect 11069 2941 11103 2975
rect 11161 2941 11195 2975
rect 11621 2941 11655 2975
rect 11713 2941 11747 2975
rect 11805 2941 11839 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 12265 2941 12299 2975
rect 12357 2941 12391 2975
rect 12541 2941 12575 2975
rect 12909 2941 12943 2975
rect 13369 2941 13403 2975
rect 13737 2941 13771 2975
rect 13829 2941 13863 2975
rect 14013 2941 14047 2975
rect 14105 2941 14139 2975
rect 14289 2941 14323 2975
rect 14381 2941 14415 2975
rect 14565 2941 14599 2975
rect 14657 2941 14691 2975
rect 14841 2941 14875 2975
rect 15853 2941 15887 2975
rect 15945 2941 15979 2975
rect 16037 2941 16071 2975
rect 16221 2941 16255 2975
rect 16313 2941 16347 2975
rect 16497 2941 16531 2975
rect 16589 2941 16623 2975
rect 16773 2941 16807 2975
rect 16865 2941 16899 2975
rect 17049 2941 17083 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 17417 2941 17451 2975
rect 17601 2941 17635 2975
rect 18521 2941 18555 2975
rect 19073 2941 19107 2975
rect 19165 2941 19199 2975
rect 19625 2941 19659 2975
rect 19717 2941 19751 2975
rect 20729 2941 20763 2975
rect 20821 2941 20855 2975
rect 21005 2941 21039 2975
rect 21097 2941 21131 2975
rect 21281 2941 21315 2975
rect 21373 2941 21407 2975
rect 21557 2941 21591 2975
rect 21649 2941 21683 2975
rect 21833 2941 21867 2975
rect 21925 2941 21959 2975
rect 22109 2941 22143 2975
rect 22201 2941 22235 2975
rect 22385 2941 22419 2975
rect 22477 2941 22511 2975
rect 22661 2941 22695 2975
rect 22753 2941 22787 2975
rect 22937 2941 22971 2975
rect 23029 2941 23063 2975
rect 23213 2941 23247 2975
rect 23305 2941 23339 2975
rect 23489 2941 23523 2975
rect 23581 2941 23615 2975
rect 23857 2941 23891 2975
rect 23949 2941 23983 2975
rect 24133 2941 24167 2975
rect 24225 2941 24259 2975
rect 24409 2941 24443 2975
rect 26525 2941 26559 2975
rect 26801 2941 26835 2975
rect 26985 2941 27019 2975
rect 27077 2941 27111 2975
rect 27169 2941 27203 2975
rect 7757 2873 7791 2907
rect 10977 2873 11011 2907
rect 19533 2873 19567 2907
rect 27261 2873 27295 2907
rect 7481 2805 7515 2839
rect 11253 2805 11287 2839
rect 13277 2805 13311 2839
rect 14933 2805 14967 2839
rect 18429 2805 18463 2839
rect 24501 2805 24535 2839
rect 11253 2601 11287 2635
rect 11805 2601 11839 2635
rect 13829 2601 13863 2635
rect 15577 2601 15611 2635
rect 15853 2601 15887 2635
rect 20729 2601 20763 2635
rect 27077 2601 27111 2635
rect 9413 2533 9447 2567
rect 10701 2533 10735 2567
rect 14197 2533 14231 2567
rect 20453 2533 20487 2567
rect 23857 2533 23891 2567
rect 7573 2465 7607 2499
rect 7665 2465 7699 2499
rect 7849 2465 7883 2499
rect 7941 2465 7975 2499
rect 8125 2465 8159 2499
rect 8217 2465 8251 2499
rect 8401 2465 8435 2499
rect 8953 2465 8987 2499
rect 9045 2465 9079 2499
rect 9321 2465 9355 2499
rect 10517 2465 10551 2499
rect 10793 2465 10827 2499
rect 11345 2465 11379 2499
rect 11437 2465 11471 2499
rect 11713 2465 11747 2499
rect 13645 2465 13679 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14381 2465 14415 2499
rect 15485 2465 15519 2499
rect 15945 2465 15979 2499
rect 16221 2465 16255 2499
rect 16313 2465 16347 2499
rect 16405 2465 16439 2499
rect 18705 2465 18739 2499
rect 18797 2465 18831 2499
rect 18889 2465 18923 2499
rect 19073 2465 19107 2499
rect 19165 2465 19199 2499
rect 19349 2465 19383 2499
rect 20545 2465 20579 2499
rect 20821 2465 20855 2499
rect 21005 2465 21039 2499
rect 21097 2465 21131 2499
rect 21281 2465 21315 2499
rect 23949 2465 23983 2499
rect 24041 2465 24075 2499
rect 24133 2465 24167 2499
rect 24317 2465 24351 2499
rect 24409 2465 24443 2499
rect 24593 2465 24627 2499
rect 24685 2465 24719 2499
rect 24869 2465 24903 2499
rect 24961 2465 24995 2499
rect 25145 2465 25179 2499
rect 25237 2465 25271 2499
rect 25421 2465 25455 2499
rect 25513 2465 25547 2499
rect 25697 2465 25731 2499
rect 25789 2465 25823 2499
rect 25973 2465 26007 2499
rect 26065 2465 26099 2499
rect 26433 2465 26467 2499
rect 26525 2465 26559 2499
rect 26709 2465 26743 2499
rect 26801 2465 26835 2499
rect 26985 2465 27019 2499
rect 8861 2397 8895 2431
rect 11529 2397 11563 2431
rect 14473 2397 14507 2431
rect 16497 2397 16531 2431
rect 19441 2397 19475 2431
rect 21373 2397 21407 2431
rect 8493 2329 8527 2363
rect 9137 2261 9171 2295
rect 10425 2261 10459 2295
rect 13553 2261 13587 2295
rect 18613 2261 18647 2295
rect 11069 2057 11103 2091
rect 11345 2057 11379 2091
rect 15577 2057 15611 2091
rect 20637 2057 20671 2091
rect 10793 1989 10827 2023
rect 8953 1921 8987 1955
rect 13921 1921 13955 1955
rect 16405 1921 16439 1955
rect 17233 1921 17267 1955
rect 19349 1921 19383 1955
rect 8769 1853 8803 1887
rect 9045 1853 9079 1887
rect 9137 1853 9171 1887
rect 9229 1853 9263 1887
rect 9413 1853 9447 1887
rect 10885 1853 10919 1887
rect 10977 1853 11011 1887
rect 11437 1853 11471 1887
rect 11621 1853 11655 1887
rect 11713 1853 11747 1887
rect 11805 1853 11839 1887
rect 12817 1853 12851 1887
rect 13001 1853 13035 1887
rect 13093 1853 13127 1887
rect 13277 1853 13311 1887
rect 13369 1853 13403 1887
rect 13553 1853 13587 1887
rect 13645 1853 13679 1887
rect 13829 1853 13863 1887
rect 15669 1853 15703 1887
rect 15853 1853 15887 1887
rect 15945 1853 15979 1887
rect 16129 1853 16163 1887
rect 16221 1853 16255 1887
rect 16313 1853 16347 1887
rect 17325 1853 17359 1887
rect 17509 1853 17543 1887
rect 17601 1853 17635 1887
rect 17693 1853 17727 1887
rect 18153 1853 18187 1887
rect 18337 1853 18371 1887
rect 18429 1853 18463 1887
rect 18797 1853 18831 1887
rect 18889 1853 18923 1887
rect 19073 1853 19107 1887
rect 19165 1853 19199 1887
rect 19257 1853 19291 1887
rect 20729 1853 20763 1887
rect 20913 1853 20947 1887
rect 21005 1853 21039 1887
rect 21189 1853 21223 1887
rect 21281 1853 21315 1887
rect 21373 1853 21407 1887
rect 9505 1785 9539 1819
rect 11897 1785 11931 1819
rect 18061 1785 18095 1819
rect 21465 1785 21499 1819
rect 8677 1717 8711 1751
rect 12725 1717 12759 1751
rect 17785 1717 17819 1751
rect 11161 1513 11195 1547
rect 15669 1513 15703 1547
rect 20637 1513 20671 1547
rect 9597 1445 9631 1479
rect 10149 1445 10183 1479
rect 11713 1445 11747 1479
rect 16497 1445 16531 1479
rect 17141 1445 17175 1479
rect 20913 1445 20947 1479
rect 21649 1445 21683 1479
rect 8677 1377 8711 1411
rect 8769 1377 8803 1411
rect 8953 1377 8987 1411
rect 9045 1377 9079 1411
rect 9413 1377 9447 1411
rect 9505 1377 9539 1411
rect 10241 1377 10275 1411
rect 10333 1377 10367 1411
rect 10425 1377 10459 1411
rect 10609 1377 10643 1411
rect 10701 1377 10735 1411
rect 11253 1377 11287 1411
rect 11437 1377 11471 1411
rect 11529 1377 11563 1411
rect 11621 1377 11655 1411
rect 13185 1377 13219 1411
rect 13277 1377 13311 1411
rect 13461 1377 13495 1411
rect 13553 1377 13587 1411
rect 13737 1377 13771 1411
rect 13829 1377 13863 1411
rect 14013 1377 14047 1411
rect 15761 1377 15795 1411
rect 16221 1377 16255 1411
rect 16313 1377 16347 1411
rect 16405 1377 16439 1411
rect 17233 1377 17267 1411
rect 17325 1377 17359 1411
rect 17417 1377 17451 1411
rect 17601 1377 17635 1411
rect 18705 1377 18739 1411
rect 18797 1377 18831 1411
rect 18981 1377 19015 1411
rect 19073 1377 19107 1411
rect 19257 1377 19291 1411
rect 19349 1377 19383 1411
rect 19533 1377 19567 1411
rect 19625 1377 19659 1411
rect 19809 1377 19843 1411
rect 20729 1377 20763 1411
rect 21005 1377 21039 1411
rect 21373 1377 21407 1411
rect 21465 1377 21499 1411
rect 21557 1377 21591 1411
rect 9321 1173 9355 1207
rect 14105 1173 14139 1207
rect 17693 1173 17727 1207
rect 19901 1173 19935 1207
rect 10425 969 10459 1003
rect 15577 969 15611 1003
rect 18797 969 18831 1003
rect 21005 969 21039 1003
rect 8861 833 8895 867
rect 9965 833 9999 867
rect 15853 833 15887 867
rect 17233 833 17267 867
rect 19809 833 19843 867
rect 8953 765 8987 799
rect 9045 765 9079 799
rect 9137 765 9171 799
rect 9321 765 9355 799
rect 9413 765 9447 799
rect 9597 765 9631 799
rect 9689 765 9723 799
rect 9873 765 9907 799
rect 10517 765 10551 799
rect 10609 765 10643 799
rect 13369 765 13403 799
rect 13737 765 13771 799
rect 13829 765 13863 799
rect 14013 765 14047 799
rect 14105 765 14139 799
rect 14289 765 14323 799
rect 14381 765 14415 799
rect 14565 765 14599 799
rect 14657 765 14691 799
rect 14841 765 14875 799
rect 14933 765 14967 799
rect 15117 765 15151 799
rect 15669 765 15703 799
rect 15761 765 15795 799
rect 17325 765 17359 799
rect 17417 765 17451 799
rect 17509 765 17543 799
rect 17693 765 17727 799
rect 17785 765 17819 799
rect 17969 765 18003 799
rect 18061 765 18095 799
rect 18245 765 18279 799
rect 18337 765 18371 799
rect 18705 765 18739 799
rect 19901 765 19935 799
rect 20085 765 20119 799
rect 20177 765 20211 799
rect 20361 765 20395 799
rect 20453 765 20487 799
rect 20637 765 20671 799
rect 20729 765 20763 799
rect 20913 765 20947 799
rect 10701 697 10735 731
rect 13277 697 13311 731
rect 15209 697 15243 731
<< metal1 >>
rect 19058 21836 19064 21888
rect 19116 21876 19122 21888
rect 26418 21876 26424 21888
rect 19116 21848 26424 21876
rect 19116 21836 19122 21848
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 552 21786 31648 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 11436 21786
rect 11488 21734 11500 21786
rect 11552 21734 11564 21786
rect 11616 21734 11628 21786
rect 11680 21734 11692 21786
rect 11744 21734 19210 21786
rect 19262 21734 19274 21786
rect 19326 21734 19338 21786
rect 19390 21734 19402 21786
rect 19454 21734 19466 21786
rect 19518 21734 26984 21786
rect 27036 21734 27048 21786
rect 27100 21734 27112 21786
rect 27164 21734 27176 21786
rect 27228 21734 27240 21786
rect 27292 21734 31648 21786
rect 552 21712 31648 21734
rect 6178 21632 6184 21684
rect 6236 21632 6242 21684
rect 6730 21632 6736 21684
rect 6788 21632 6794 21684
rect 7282 21632 7288 21684
rect 7340 21632 7346 21684
rect 7834 21632 7840 21684
rect 7892 21632 7898 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 8938 21632 8944 21684
rect 8996 21632 9002 21684
rect 9490 21632 9496 21684
rect 9548 21632 9554 21684
rect 10042 21632 10048 21684
rect 10100 21632 10106 21684
rect 10594 21632 10600 21684
rect 10652 21632 10658 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11701 21675 11759 21681
rect 11701 21641 11713 21675
rect 11747 21672 11759 21675
rect 11790 21672 11796 21684
rect 11747 21644 11796 21672
rect 11747 21641 11759 21644
rect 11701 21635 11759 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 13538 21632 13544 21684
rect 13596 21632 13602 21684
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 14458 21632 14464 21684
rect 14516 21632 14522 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 15381 21675 15439 21681
rect 15381 21672 15393 21675
rect 15252 21644 15393 21672
rect 15252 21632 15258 21644
rect 15381 21641 15393 21644
rect 15427 21641 15439 21675
rect 15381 21635 15439 21641
rect 15654 21632 15660 21684
rect 15712 21632 15718 21684
rect 16114 21632 16120 21684
rect 16172 21632 16178 21684
rect 16758 21632 16764 21684
rect 16816 21632 16822 21684
rect 16942 21632 16948 21684
rect 17000 21632 17006 21684
rect 17586 21632 17592 21684
rect 17644 21632 17650 21684
rect 18322 21632 18328 21684
rect 18380 21632 18386 21684
rect 19889 21675 19947 21681
rect 19889 21641 19901 21675
rect 19935 21672 19947 21675
rect 19935 21644 23152 21672
rect 19935 21641 19947 21644
rect 19889 21635 19947 21641
rect 19058 21604 19064 21616
rect 15580 21576 19064 21604
rect 15580 21477 15608 21576
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 23124 21613 23152 21644
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 24673 21675 24731 21681
rect 24673 21672 24685 21675
rect 23256 21644 24685 21672
rect 23256 21632 23262 21644
rect 24673 21641 24685 21644
rect 24719 21641 24731 21675
rect 24673 21635 24731 21641
rect 24857 21675 24915 21681
rect 24857 21641 24869 21675
rect 24903 21672 24915 21675
rect 26050 21672 26056 21684
rect 24903 21644 26056 21672
rect 24903 21641 24915 21644
rect 24857 21635 24915 21641
rect 26050 21632 26056 21644
rect 26108 21632 26114 21684
rect 26418 21632 26424 21684
rect 26476 21632 26482 21684
rect 27065 21675 27123 21681
rect 27065 21672 27077 21675
rect 26620 21644 27077 21672
rect 19429 21607 19487 21613
rect 19429 21604 19441 21607
rect 19392 21576 19441 21604
rect 19392 21564 19398 21576
rect 19429 21573 19441 21576
rect 19475 21573 19487 21607
rect 19429 21567 19487 21573
rect 20533 21607 20591 21613
rect 20533 21573 20545 21607
rect 20579 21604 20591 21607
rect 22097 21607 22155 21613
rect 20579 21576 22048 21604
rect 20579 21573 20591 21576
rect 20533 21567 20591 21573
rect 19794 21536 19800 21548
rect 19628 21508 19800 21536
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21437 15623 21471
rect 15565 21431 15623 21437
rect 16574 21428 16580 21480
rect 16632 21428 16638 21480
rect 17402 21428 17408 21480
rect 17460 21428 17466 21480
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21468 18567 21471
rect 18874 21468 18880 21480
rect 18555 21440 18880 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 19628 21477 19656 21508
rect 19794 21496 19800 21508
rect 19852 21536 19858 21548
rect 20165 21539 20223 21545
rect 20165 21536 20177 21539
rect 19852 21508 20177 21536
rect 19852 21496 19858 21508
rect 20165 21505 20177 21508
rect 20211 21505 20223 21539
rect 20165 21499 20223 21505
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 22020 21536 22048 21576
rect 22097 21573 22109 21607
rect 22143 21604 22155 21607
rect 22189 21607 22247 21613
rect 22189 21604 22201 21607
rect 22143 21576 22201 21604
rect 22143 21573 22155 21576
rect 22097 21567 22155 21573
rect 22189 21573 22201 21576
rect 22235 21573 22247 21607
rect 22189 21567 22247 21573
rect 23109 21607 23167 21613
rect 23109 21573 23121 21607
rect 23155 21573 23167 21607
rect 23109 21567 23167 21573
rect 24949 21607 25007 21613
rect 24949 21573 24961 21607
rect 24995 21573 25007 21607
rect 26620 21604 26648 21644
rect 27065 21641 27077 21644
rect 27111 21641 27123 21675
rect 27065 21635 27123 21641
rect 24949 21567 25007 21573
rect 25332 21576 26648 21604
rect 26973 21607 27031 21613
rect 24964 21536 24992 21567
rect 20772 21508 21312 21536
rect 22020 21508 23336 21536
rect 20772 21496 20778 21508
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21437 19671 21471
rect 19613 21431 19671 21437
rect 19702 21428 19708 21480
rect 19760 21428 19766 21480
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 20272 21400 20300 21431
rect 20346 21428 20352 21480
rect 20404 21428 20410 21480
rect 20809 21471 20867 21477
rect 20809 21437 20821 21471
rect 20855 21468 20867 21471
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20855 21440 21005 21468
rect 20855 21437 20867 21440
rect 20809 21431 20867 21437
rect 20993 21437 21005 21440
rect 21039 21437 21051 21471
rect 20993 21431 21051 21437
rect 21082 21428 21088 21480
rect 21140 21428 21146 21480
rect 21284 21477 21312 21508
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21437 21327 21471
rect 21269 21431 21327 21437
rect 21545 21471 21603 21477
rect 21545 21437 21557 21471
rect 21591 21468 21603 21471
rect 21591 21440 22048 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 20717 21403 20775 21409
rect 20717 21400 20729 21403
rect 20272 21372 20729 21400
rect 20717 21369 20729 21372
rect 20763 21369 20775 21403
rect 21821 21403 21879 21409
rect 21821 21400 21833 21403
rect 20717 21363 20775 21369
rect 21468 21372 21833 21400
rect 21468 21341 21496 21372
rect 21821 21369 21833 21372
rect 21867 21369 21879 21403
rect 22020 21400 22048 21440
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22373 21471 22431 21477
rect 22373 21468 22385 21471
rect 22152 21440 22385 21468
rect 22152 21428 22158 21440
rect 22373 21437 22385 21440
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 22646 21428 22652 21480
rect 22704 21428 22710 21480
rect 22738 21428 22744 21480
rect 22796 21428 22802 21480
rect 23198 21468 23204 21480
rect 23124 21440 23204 21468
rect 23124 21400 23152 21440
rect 23198 21428 23204 21440
rect 23256 21428 23262 21480
rect 23308 21477 23336 21508
rect 24044 21508 24992 21536
rect 24044 21477 24072 21508
rect 23293 21471 23351 21477
rect 23293 21437 23305 21471
rect 23339 21437 23351 21471
rect 23293 21431 23351 21437
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21468 23719 21471
rect 24029 21471 24087 21477
rect 23707 21440 23980 21468
rect 23707 21437 23719 21440
rect 23661 21431 23719 21437
rect 22020 21372 23152 21400
rect 23216 21372 23796 21400
rect 21821 21363 21879 21369
rect 21453 21335 21511 21341
rect 21453 21301 21465 21335
rect 21499 21301 21511 21335
rect 21453 21295 21511 21301
rect 21726 21292 21732 21344
rect 21784 21292 21790 21344
rect 21913 21335 21971 21341
rect 21913 21301 21925 21335
rect 21959 21332 21971 21335
rect 22465 21335 22523 21341
rect 22465 21332 22477 21335
rect 21959 21304 22477 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22465 21301 22477 21304
rect 22511 21301 22523 21335
rect 22465 21295 22523 21301
rect 22925 21335 22983 21341
rect 22925 21301 22937 21335
rect 22971 21332 22983 21335
rect 23216 21332 23244 21372
rect 22971 21304 23244 21332
rect 22971 21301 22983 21304
rect 22925 21295 22983 21301
rect 23290 21292 23296 21344
rect 23348 21332 23354 21344
rect 23385 21335 23443 21341
rect 23385 21332 23397 21335
rect 23348 21304 23397 21332
rect 23348 21292 23354 21304
rect 23385 21301 23397 21304
rect 23431 21301 23443 21335
rect 23385 21295 23443 21301
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23658 21332 23664 21344
rect 23523 21304 23664 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 23768 21332 23796 21372
rect 23842 21360 23848 21412
rect 23900 21360 23906 21412
rect 23952 21400 23980 21440
rect 24029 21437 24041 21471
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24912 21440 25145 21468
rect 24912 21428 24918 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25332 21468 25360 21576
rect 26973 21573 26985 21607
rect 27019 21604 27031 21607
rect 27341 21607 27399 21613
rect 27341 21604 27353 21607
rect 27019 21576 27353 21604
rect 27019 21573 27031 21576
rect 26973 21567 27031 21573
rect 27341 21573 27353 21576
rect 27387 21573 27399 21607
rect 27341 21567 27399 21573
rect 28166 21564 28172 21616
rect 28224 21604 28230 21616
rect 29549 21607 29607 21613
rect 29549 21604 29561 21607
rect 28224 21576 29561 21604
rect 28224 21564 28230 21576
rect 29549 21573 29561 21576
rect 29595 21573 29607 21607
rect 29549 21567 29607 21573
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21536 25467 21539
rect 29089 21539 29147 21545
rect 29089 21536 29101 21539
rect 25455 21508 26740 21536
rect 25455 21505 25467 21508
rect 25409 21499 25467 21505
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 25332 21440 25789 21468
rect 25133 21431 25191 21437
rect 25777 21437 25789 21440
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21468 26295 21471
rect 26326 21468 26332 21480
rect 26283 21440 26332 21468
rect 26283 21437 26295 21440
rect 26237 21431 26295 21437
rect 26326 21428 26332 21440
rect 26384 21428 26390 21480
rect 26712 21477 26740 21508
rect 28368 21508 29101 21536
rect 26697 21471 26755 21477
rect 26697 21437 26709 21471
rect 26743 21437 26755 21471
rect 26697 21431 26755 21437
rect 27246 21428 27252 21480
rect 27304 21428 27310 21480
rect 27522 21428 27528 21480
rect 27580 21428 27586 21480
rect 28368 21477 28396 21508
rect 29089 21505 29101 21508
rect 29135 21505 29147 21539
rect 29089 21499 29147 21505
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21468 27859 21471
rect 27985 21471 28043 21477
rect 27985 21468 27997 21471
rect 27847 21440 27997 21468
rect 27847 21437 27859 21440
rect 27801 21431 27859 21437
rect 27985 21437 27997 21440
rect 28031 21437 28043 21471
rect 27985 21431 28043 21437
rect 28077 21471 28135 21477
rect 28077 21437 28089 21471
rect 28123 21468 28135 21471
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 28123 21440 28273 21468
rect 28123 21437 28135 21440
rect 28077 21431 28135 21437
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21437 28411 21471
rect 28353 21431 28411 21437
rect 28626 21428 28632 21480
rect 28684 21428 28690 21480
rect 28994 21428 29000 21480
rect 29052 21428 29058 21480
rect 29454 21428 29460 21480
rect 29512 21428 29518 21480
rect 29730 21428 29736 21480
rect 29788 21428 29794 21480
rect 24489 21403 24547 21409
rect 24489 21400 24501 21403
rect 23952 21372 24501 21400
rect 24489 21369 24501 21372
rect 24535 21369 24547 21403
rect 24489 21363 24547 21369
rect 25593 21403 25651 21409
rect 25593 21369 25605 21403
rect 25639 21400 25651 21403
rect 25639 21372 25912 21400
rect 25639 21369 25651 21372
rect 25593 21363 25651 21369
rect 24121 21335 24179 21341
rect 24121 21332 24133 21335
rect 23768 21304 24133 21332
rect 24121 21301 24133 21304
rect 24167 21301 24179 21335
rect 24121 21295 24179 21301
rect 24210 21292 24216 21344
rect 24268 21292 24274 21344
rect 24397 21335 24455 21341
rect 24397 21301 24409 21335
rect 24443 21332 24455 21335
rect 24689 21335 24747 21341
rect 24689 21332 24701 21335
rect 24443 21304 24701 21332
rect 24443 21301 24455 21304
rect 24397 21295 24455 21301
rect 24689 21301 24701 21304
rect 24735 21301 24747 21335
rect 24689 21295 24747 21301
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 25884 21332 25912 21372
rect 25958 21360 25964 21412
rect 26016 21360 26022 21412
rect 26068 21400 26096 21428
rect 26605 21403 26663 21409
rect 26605 21400 26617 21403
rect 26068 21372 26617 21400
rect 26605 21369 26617 21372
rect 26651 21369 26663 21403
rect 26605 21363 26663 21369
rect 26789 21403 26847 21409
rect 26789 21369 26801 21403
rect 26835 21400 26847 21403
rect 26835 21372 28488 21400
rect 26835 21369 26847 21372
rect 26789 21363 26847 21369
rect 26053 21335 26111 21341
rect 26053 21332 26065 21335
rect 25884 21304 26065 21332
rect 26053 21301 26065 21304
rect 26099 21301 26111 21335
rect 26053 21295 26111 21301
rect 27709 21335 27767 21341
rect 27709 21301 27721 21335
rect 27755 21332 27767 21335
rect 28074 21332 28080 21344
rect 27755 21304 28080 21332
rect 27755 21301 27767 21304
rect 27709 21295 27767 21301
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 28460 21341 28488 21372
rect 28445 21335 28503 21341
rect 28445 21301 28457 21335
rect 28491 21301 28503 21335
rect 28445 21295 28503 21301
rect 29270 21292 29276 21344
rect 29328 21332 29334 21344
rect 29365 21335 29423 21341
rect 29365 21332 29377 21335
rect 29328 21304 29377 21332
rect 29328 21292 29334 21304
rect 29365 21301 29377 21304
rect 29411 21301 29423 21335
rect 29365 21295 29423 21301
rect 552 21242 31648 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 12096 21242
rect 12148 21190 12160 21242
rect 12212 21190 12224 21242
rect 12276 21190 12288 21242
rect 12340 21190 12352 21242
rect 12404 21190 19870 21242
rect 19922 21190 19934 21242
rect 19986 21190 19998 21242
rect 20050 21190 20062 21242
rect 20114 21190 20126 21242
rect 20178 21190 27644 21242
rect 27696 21190 27708 21242
rect 27760 21190 27772 21242
rect 27824 21190 27836 21242
rect 27888 21190 27900 21242
rect 27952 21190 31648 21242
rect 552 21168 31648 21190
rect 15381 21131 15439 21137
rect 15381 21097 15393 21131
rect 15427 21128 15439 21131
rect 16574 21128 16580 21140
rect 15427 21100 16580 21128
rect 15427 21097 15439 21100
rect 15381 21091 15439 21097
rect 15396 21060 15424 21091
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 21082 21088 21088 21140
rect 21140 21128 21146 21140
rect 21361 21131 21419 21137
rect 21361 21128 21373 21131
rect 21140 21100 21373 21128
rect 21140 21088 21146 21100
rect 21361 21097 21373 21100
rect 21407 21097 21419 21131
rect 21361 21091 21419 21097
rect 21726 21088 21732 21140
rect 21784 21088 21790 21140
rect 23661 21131 23719 21137
rect 23661 21097 23673 21131
rect 23707 21097 23719 21131
rect 23661 21091 23719 21097
rect 17589 21063 17647 21069
rect 17589 21060 17601 21063
rect 15212 21032 15424 21060
rect 17420 21032 17601 21060
rect 12342 20952 12348 21004
rect 12400 20952 12406 21004
rect 15212 21001 15240 21032
rect 17420 21004 17448 21032
rect 17589 21029 17601 21032
rect 17635 21029 17647 21063
rect 17589 21023 17647 21029
rect 19794 21020 19800 21072
rect 19852 21060 19858 21072
rect 23676 21060 23704 21091
rect 23842 21088 23848 21140
rect 23900 21088 23906 21140
rect 25133 21131 25191 21137
rect 25133 21097 25145 21131
rect 25179 21128 25191 21131
rect 25682 21128 25688 21140
rect 25179 21100 25688 21128
rect 25179 21097 25191 21100
rect 25133 21091 25191 21097
rect 25682 21088 25688 21100
rect 25740 21088 25746 21140
rect 25958 21088 25964 21140
rect 26016 21128 26022 21140
rect 26053 21131 26111 21137
rect 26053 21128 26065 21131
rect 26016 21100 26065 21128
rect 26016 21088 26022 21100
rect 26053 21097 26065 21100
rect 26099 21097 26111 21131
rect 28166 21128 28172 21140
rect 26053 21091 26111 21097
rect 26206 21100 28172 21128
rect 24210 21060 24216 21072
rect 19852 21032 20116 21060
rect 23676 21032 24216 21060
rect 19852 21020 19858 21032
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 12621 20995 12679 21001
rect 12621 20992 12633 20995
rect 12483 20964 12633 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 12621 20961 12633 20964
rect 12667 20961 12679 20995
rect 12621 20955 12679 20961
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12759 20964 12909 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 12989 20995 13047 21001
rect 12989 20961 13001 20995
rect 13035 20992 13047 20995
rect 13173 20995 13231 21001
rect 13173 20992 13185 20995
rect 13035 20964 13185 20992
rect 13035 20961 13047 20964
rect 12989 20955 13047 20961
rect 13173 20961 13185 20964
rect 13219 20961 13231 20995
rect 13173 20955 13231 20961
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 13541 20995 13599 21001
rect 13541 20992 13553 20995
rect 13311 20964 13553 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 13541 20961 13553 20964
rect 13587 20961 13599 20995
rect 13541 20955 13599 20961
rect 13633 20995 13691 21001
rect 13633 20961 13645 20995
rect 13679 20992 13691 20995
rect 13909 20995 13967 21001
rect 13909 20992 13921 20995
rect 13679 20964 13921 20992
rect 13679 20961 13691 20964
rect 13633 20955 13691 20961
rect 13909 20961 13921 20964
rect 13955 20961 13967 20995
rect 13909 20955 13967 20961
rect 14001 20995 14059 21001
rect 14001 20961 14013 20995
rect 14047 20992 14059 20995
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 14047 20964 14289 20992
rect 14047 20961 14059 20964
rect 14001 20955 14059 20961
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 14967 20964 15117 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20961 15255 20995
rect 15197 20955 15255 20961
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20961 15347 20995
rect 15289 20955 15347 20961
rect 16577 20995 16635 21001
rect 16577 20961 16589 20995
rect 16623 20992 16635 20995
rect 16761 20995 16819 21001
rect 16761 20992 16773 20995
rect 16623 20964 16773 20992
rect 16623 20961 16635 20964
rect 16577 20955 16635 20961
rect 16761 20961 16773 20964
rect 16807 20961 16819 20995
rect 16761 20955 16819 20961
rect 16853 20995 16911 21001
rect 16853 20961 16865 20995
rect 16899 20992 16911 20995
rect 17037 20995 17095 21001
rect 17037 20992 17049 20995
rect 16899 20964 17049 20992
rect 16899 20961 16911 20964
rect 16853 20955 16911 20961
rect 17037 20961 17049 20964
rect 17083 20961 17095 20995
rect 17037 20955 17095 20961
rect 17129 20995 17187 21001
rect 17129 20961 17141 20995
rect 17175 20992 17187 20995
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 17175 20964 17325 20992
rect 17175 20961 17187 20964
rect 17129 20955 17187 20961
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 15304 20924 15332 20955
rect 17402 20952 17408 21004
rect 17460 20952 17466 21004
rect 17494 20952 17500 21004
rect 17552 20952 17558 21004
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20992 18659 20995
rect 18785 20995 18843 21001
rect 18785 20992 18797 20995
rect 18647 20964 18797 20992
rect 18647 20961 18659 20964
rect 18601 20955 18659 20961
rect 18785 20961 18797 20964
rect 18831 20961 18843 20995
rect 18785 20955 18843 20961
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 19061 20995 19119 21001
rect 19061 20992 19073 20995
rect 18932 20964 19073 20992
rect 18932 20952 18938 20964
rect 19061 20961 19073 20964
rect 19107 20961 19119 20995
rect 19061 20955 19119 20961
rect 19153 20995 19211 21001
rect 19153 20961 19165 20995
rect 19199 20992 19211 20995
rect 19337 20995 19395 21001
rect 19337 20992 19349 20995
rect 19199 20964 19349 20992
rect 19199 20961 19211 20964
rect 19153 20955 19211 20961
rect 19337 20961 19349 20964
rect 19383 20961 19395 20995
rect 19337 20955 19395 20961
rect 19429 20995 19487 21001
rect 19429 20961 19441 20995
rect 19475 20992 19487 20995
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19475 20964 19625 20992
rect 19475 20961 19487 20964
rect 19429 20955 19487 20961
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 19613 20955 19671 20961
rect 19705 20995 19763 21001
rect 19705 20961 19717 20995
rect 19751 20992 19763 20995
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19751 20964 19901 20992
rect 19751 20961 19763 20964
rect 19705 20955 19763 20961
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 19978 20952 19984 21004
rect 20036 20952 20042 21004
rect 20088 21001 20116 21032
rect 24210 21020 24216 21032
rect 24268 21020 24274 21072
rect 26206 21060 26234 21100
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 28445 21131 28503 21137
rect 28445 21097 28457 21131
rect 28491 21128 28503 21131
rect 28994 21128 29000 21140
rect 28491 21100 29000 21128
rect 28491 21097 28503 21100
rect 28445 21091 28503 21097
rect 28994 21088 29000 21100
rect 29052 21088 29058 21140
rect 29454 21088 29460 21140
rect 29512 21128 29518 21140
rect 29917 21131 29975 21137
rect 29917 21128 29929 21131
rect 29512 21100 29929 21128
rect 29512 21088 29518 21100
rect 29917 21097 29929 21100
rect 29963 21097 29975 21131
rect 29917 21091 29975 21097
rect 27985 21063 28043 21069
rect 27985 21060 27997 21063
rect 24872 21032 26234 21060
rect 27816 21032 27997 21060
rect 20073 20995 20131 21001
rect 20073 20961 20085 20995
rect 20119 20961 20131 20995
rect 20073 20955 20131 20961
rect 20165 20995 20223 21001
rect 20165 20961 20177 20995
rect 20211 20992 20223 20995
rect 20349 20995 20407 21001
rect 20349 20992 20361 20995
rect 20211 20964 20361 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 20349 20961 20361 20964
rect 20395 20961 20407 20995
rect 20349 20955 20407 20961
rect 20441 20995 20499 21001
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 20487 20964 20637 20992
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 20625 20955 20683 20961
rect 21453 20995 21511 21001
rect 21453 20961 21465 20995
rect 21499 20961 21511 20995
rect 21453 20955 21511 20961
rect 14415 20896 15332 20924
rect 21468 20924 21496 20955
rect 21542 20952 21548 21004
rect 21600 20952 21606 21004
rect 22005 20995 22063 21001
rect 22005 20961 22017 20995
rect 22051 20992 22063 20995
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 22051 20964 22201 20992
rect 22051 20961 22063 20964
rect 22005 20955 22063 20961
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 22281 20995 22339 21001
rect 22281 20961 22293 20995
rect 22327 20992 22339 20995
rect 22465 20995 22523 21001
rect 22465 20992 22477 20995
rect 22327 20964 22477 20992
rect 22327 20961 22339 20964
rect 22281 20955 22339 20961
rect 22465 20961 22477 20964
rect 22511 20961 22523 20995
rect 22465 20955 22523 20961
rect 22557 20995 22615 21001
rect 22557 20961 22569 20995
rect 22603 20992 22615 20995
rect 22741 20995 22799 21001
rect 22741 20992 22753 20995
rect 22603 20964 22753 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 22741 20961 22753 20964
rect 22787 20961 22799 20995
rect 22741 20955 22799 20961
rect 22833 20995 22891 21001
rect 22833 20961 22845 20995
rect 22879 20992 22891 20995
rect 23017 20995 23075 21001
rect 23017 20992 23029 20995
rect 22879 20964 23029 20992
rect 22879 20961 22891 20964
rect 22833 20955 22891 20961
rect 23017 20961 23029 20964
rect 23063 20961 23075 20995
rect 23017 20955 23075 20961
rect 23109 20995 23167 21001
rect 23109 20961 23121 20995
rect 23155 20992 23167 20995
rect 23293 20995 23351 21001
rect 23293 20992 23305 20995
rect 23155 20964 23305 20992
rect 23155 20961 23167 20964
rect 23109 20955 23167 20961
rect 23293 20961 23305 20964
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23382 20952 23388 21004
rect 23440 20952 23446 21004
rect 23474 20952 23480 21004
rect 23532 20952 23538 21004
rect 24026 20952 24032 21004
rect 24084 20952 24090 21004
rect 21913 20927 21971 20933
rect 21913 20924 21925 20927
rect 21468 20896 21925 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 21913 20893 21925 20896
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 23658 20884 23664 20936
rect 23716 20924 23722 20936
rect 24872 20924 24900 21032
rect 24946 20952 24952 21004
rect 25004 20952 25010 21004
rect 26234 20952 26240 21004
rect 26292 20952 26298 21004
rect 27816 21001 27844 21032
rect 27985 21029 27997 21032
rect 28031 21029 28043 21063
rect 29365 21063 29423 21069
rect 29365 21060 29377 21063
rect 27985 21023 28043 21029
rect 28552 21032 29377 21060
rect 26973 20995 27031 21001
rect 26973 20961 26985 20995
rect 27019 20992 27031 20995
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 27019 20964 27169 20992
rect 27019 20961 27031 20964
rect 26973 20955 27031 20961
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 27249 20995 27307 21001
rect 27249 20961 27261 20995
rect 27295 20992 27307 20995
rect 27433 20995 27491 21001
rect 27433 20992 27445 20995
rect 27295 20964 27445 20992
rect 27295 20961 27307 20964
rect 27249 20955 27307 20961
rect 27433 20961 27445 20964
rect 27479 20961 27491 20995
rect 27433 20955 27491 20961
rect 27525 20995 27583 21001
rect 27525 20961 27537 20995
rect 27571 20992 27583 20995
rect 27709 20995 27767 21001
rect 27709 20992 27721 20995
rect 27571 20964 27721 20992
rect 27571 20961 27583 20964
rect 27525 20955 27583 20961
rect 27709 20961 27721 20964
rect 27755 20961 27767 20995
rect 27709 20955 27767 20961
rect 27801 20995 27859 21001
rect 27801 20961 27813 20995
rect 27847 20961 27859 20995
rect 27801 20955 27859 20961
rect 27893 20995 27951 21001
rect 27893 20961 27905 20995
rect 27939 20992 27951 20995
rect 28074 20992 28080 21004
rect 27939 20964 28080 20992
rect 27939 20961 27951 20964
rect 27893 20955 27951 20961
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 28552 21001 28580 21032
rect 29365 21029 29377 21032
rect 29411 21029 29423 21063
rect 29365 21023 29423 21029
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20961 28595 20995
rect 28537 20955 28595 20961
rect 28810 20952 28816 21004
rect 28868 20952 28874 21004
rect 29178 20952 29184 21004
rect 29236 20952 29242 21004
rect 29270 20952 29276 21004
rect 29328 20952 29334 21004
rect 29549 20995 29607 21001
rect 29549 20961 29561 20995
rect 29595 20961 29607 20995
rect 29549 20955 29607 20961
rect 29641 20995 29699 21001
rect 29641 20961 29653 20995
rect 29687 20992 29699 20995
rect 29825 20995 29883 21001
rect 29825 20992 29837 20995
rect 29687 20964 29837 20992
rect 29687 20961 29699 20964
rect 29641 20955 29699 20961
rect 29825 20961 29837 20964
rect 29871 20961 29883 20995
rect 29825 20955 29883 20961
rect 23716 20896 24900 20924
rect 29089 20927 29147 20933
rect 23716 20884 23722 20896
rect 29089 20893 29101 20927
rect 29135 20924 29147 20927
rect 29564 20924 29592 20955
rect 29135 20896 29592 20924
rect 29135 20893 29147 20896
rect 29089 20887 29147 20893
rect 23290 20816 23296 20868
rect 23348 20856 23354 20868
rect 28629 20859 28687 20865
rect 28629 20856 28641 20859
rect 23348 20828 28641 20856
rect 23348 20816 23354 20828
rect 28629 20825 28641 20828
rect 28675 20825 28687 20859
rect 28629 20819 28687 20825
rect 14829 20791 14887 20797
rect 14829 20757 14841 20791
rect 14875 20788 14887 20791
rect 15010 20788 15016 20800
rect 14875 20760 15016 20788
rect 14875 20757 14887 20760
rect 14829 20751 14887 20757
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 16482 20748 16488 20800
rect 16540 20748 16546 20800
rect 18506 20748 18512 20800
rect 18564 20748 18570 20800
rect 20717 20791 20775 20797
rect 20717 20757 20729 20791
rect 20763 20788 20775 20791
rect 20806 20788 20812 20800
rect 20763 20760 20812 20788
rect 20763 20757 20775 20760
rect 20717 20751 20775 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 26881 20791 26939 20797
rect 26881 20757 26893 20791
rect 26927 20788 26939 20791
rect 27430 20788 27436 20800
rect 26927 20760 27436 20788
rect 26927 20757 26939 20760
rect 26881 20751 26939 20757
rect 27430 20748 27436 20760
rect 27488 20748 27494 20800
rect 552 20698 31648 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 11436 20698
rect 11488 20646 11500 20698
rect 11552 20646 11564 20698
rect 11616 20646 11628 20698
rect 11680 20646 11692 20698
rect 11744 20646 19210 20698
rect 19262 20646 19274 20698
rect 19326 20646 19338 20698
rect 19390 20646 19402 20698
rect 19454 20646 19466 20698
rect 19518 20646 26984 20698
rect 27036 20646 27048 20698
rect 27100 20646 27112 20698
rect 27164 20646 27176 20698
rect 27228 20646 27240 20698
rect 27292 20646 31648 20698
rect 552 20624 31648 20646
rect 12342 20544 12348 20596
rect 12400 20544 12406 20596
rect 17494 20544 17500 20596
rect 17552 20544 17558 20596
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 19978 20584 19984 20596
rect 19935 20556 19984 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 23293 20587 23351 20593
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 23382 20584 23388 20596
rect 23339 20556 23388 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 29178 20544 29184 20596
rect 29236 20584 29242 20596
rect 29641 20587 29699 20593
rect 29641 20584 29653 20587
rect 29236 20556 29653 20584
rect 29236 20544 29242 20556
rect 29641 20553 29653 20556
rect 29687 20553 29699 20587
rect 29641 20547 29699 20553
rect 8481 20451 8539 20457
rect 8481 20448 8493 20451
rect 8128 20420 8493 20448
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 1581 20383 1639 20389
rect 1581 20380 1593 20383
rect 1452 20352 1593 20380
rect 1452 20340 1458 20352
rect 1581 20349 1593 20352
rect 1627 20349 1639 20383
rect 1581 20343 1639 20349
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 1118 20272 1124 20324
rect 1176 20312 1182 20324
rect 1872 20312 1900 20343
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3789 20383 3847 20389
rect 3789 20380 3801 20383
rect 3384 20352 3801 20380
rect 3384 20340 3390 20352
rect 3789 20349 3801 20352
rect 3835 20349 3847 20383
rect 3789 20343 3847 20349
rect 6454 20340 6460 20392
rect 6512 20340 6518 20392
rect 8128 20389 8156 20420
rect 8481 20417 8493 20420
rect 8527 20417 8539 20451
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 8481 20411 8539 20417
rect 12176 20420 12633 20448
rect 6549 20383 6607 20389
rect 6549 20349 6561 20383
rect 6595 20380 6607 20383
rect 6733 20383 6791 20389
rect 6733 20380 6745 20383
rect 6595 20352 6745 20380
rect 6595 20349 6607 20352
rect 6549 20343 6607 20349
rect 6733 20349 6745 20352
rect 6779 20349 6791 20383
rect 6733 20343 6791 20349
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 6871 20352 7021 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20380 7159 20383
rect 7285 20383 7343 20389
rect 7285 20380 7297 20383
rect 7147 20352 7297 20380
rect 7147 20349 7159 20352
rect 7101 20343 7159 20349
rect 7285 20349 7297 20352
rect 7331 20349 7343 20383
rect 7285 20343 7343 20349
rect 7377 20383 7435 20389
rect 7377 20349 7389 20383
rect 7423 20380 7435 20383
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 7423 20352 7573 20380
rect 7423 20349 7435 20352
rect 7377 20343 7435 20349
rect 7561 20349 7573 20352
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20349 8171 20383
rect 8113 20343 8171 20349
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 1176 20284 1900 20312
rect 7653 20315 7711 20321
rect 1176 20272 1182 20284
rect 7653 20281 7665 20315
rect 7699 20312 7711 20315
rect 8404 20312 8432 20343
rect 11238 20340 11244 20392
rect 11296 20340 11302 20392
rect 12176 20389 12204 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 15105 20451 15163 20457
rect 15105 20448 15117 20451
rect 12621 20411 12679 20417
rect 14660 20420 15117 20448
rect 14660 20389 14688 20420
rect 15105 20417 15117 20420
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 18417 20451 18475 20457
rect 17267 20420 17448 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 11333 20383 11391 20389
rect 11333 20349 11345 20383
rect 11379 20349 11391 20383
rect 11333 20343 11391 20349
rect 11425 20383 11483 20389
rect 11425 20349 11437 20383
rect 11471 20380 11483 20383
rect 11609 20383 11667 20389
rect 11609 20380 11621 20383
rect 11471 20352 11621 20380
rect 11471 20349 11483 20352
rect 11425 20343 11483 20349
rect 11609 20349 11621 20352
rect 11655 20349 11667 20383
rect 11609 20343 11667 20349
rect 12161 20383 12219 20389
rect 12161 20349 12173 20383
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20349 14703 20383
rect 14645 20343 14703 20349
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20349 14795 20383
rect 14737 20343 14795 20349
rect 7699 20284 8432 20312
rect 11149 20315 11207 20321
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 11149 20281 11161 20315
rect 11195 20312 11207 20315
rect 11348 20312 11376 20343
rect 11195 20284 11376 20312
rect 12069 20315 12127 20321
rect 11195 20281 11207 20284
rect 11149 20275 11207 20281
rect 12069 20281 12081 20315
rect 12115 20312 12127 20315
rect 12268 20312 12296 20343
rect 12115 20284 12296 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 1210 20204 1216 20256
rect 1268 20244 1274 20256
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1268 20216 1685 20244
rect 1268 20204 1274 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 1673 20207 1731 20213
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 1949 20247 2007 20253
rect 1949 20244 1961 20247
rect 1820 20216 1961 20244
rect 1820 20204 1826 20216
rect 1949 20213 1961 20216
rect 1995 20213 2007 20247
rect 1949 20207 2007 20213
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 3881 20247 3939 20253
rect 3881 20244 3893 20247
rect 3752 20216 3893 20244
rect 3752 20204 3758 20216
rect 3881 20213 3893 20216
rect 3927 20213 3939 20247
rect 3881 20207 3939 20213
rect 8021 20247 8079 20253
rect 8021 20213 8033 20247
rect 8067 20244 8079 20247
rect 8754 20244 8760 20256
rect 8067 20216 8760 20244
rect 8067 20213 8079 20216
rect 8021 20207 8079 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12544 20244 12572 20343
rect 14553 20315 14611 20321
rect 14553 20281 14565 20315
rect 14599 20312 14611 20315
rect 14752 20312 14780 20343
rect 15010 20340 15016 20392
rect 15068 20340 15074 20392
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20380 16267 20383
rect 16393 20383 16451 20389
rect 16393 20380 16405 20383
rect 16255 20352 16405 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 16393 20349 16405 20352
rect 16439 20349 16451 20383
rect 16393 20343 16451 20349
rect 16482 20340 16488 20392
rect 16540 20340 16546 20392
rect 17310 20340 17316 20392
rect 17368 20340 17374 20392
rect 17420 20389 17448 20420
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 19613 20451 19671 20457
rect 18463 20420 18736 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 18506 20340 18512 20392
rect 18564 20340 18570 20392
rect 18708 20389 18736 20420
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 24489 20451 24547 20457
rect 24489 20448 24501 20451
rect 19659 20420 19840 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20349 18751 20383
rect 18693 20343 18751 20349
rect 19702 20340 19708 20392
rect 19760 20340 19766 20392
rect 19812 20389 19840 20420
rect 24320 20420 24501 20448
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 20806 20340 20812 20392
rect 20864 20340 20870 20392
rect 24320 20389 24348 20420
rect 24489 20417 24501 20420
rect 24535 20417 24547 20451
rect 24489 20411 24547 20417
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20380 20959 20383
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 20947 20352 21097 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21085 20349 21097 20352
rect 21131 20349 21143 20383
rect 21085 20343 21143 20349
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 21223 20352 21373 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 23385 20383 23443 20389
rect 23385 20349 23397 20383
rect 23431 20380 23443 20383
rect 23569 20383 23627 20389
rect 23569 20380 23581 20383
rect 23431 20352 23581 20380
rect 23431 20349 23443 20352
rect 23385 20343 23443 20349
rect 23569 20349 23581 20352
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 23661 20383 23719 20389
rect 23661 20349 23673 20383
rect 23707 20380 23719 20383
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23707 20352 23949 20380
rect 23707 20349 23719 20352
rect 23661 20343 23719 20349
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 24029 20383 24087 20389
rect 24029 20349 24041 20383
rect 24075 20380 24087 20383
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 24075 20352 24225 20380
rect 24075 20349 24087 20352
rect 24029 20343 24087 20349
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 24305 20383 24363 20389
rect 24305 20349 24317 20383
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 24394 20340 24400 20392
rect 24452 20340 24458 20392
rect 26789 20383 26847 20389
rect 26789 20349 26801 20383
rect 26835 20380 26847 20383
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26835 20352 26985 20380
rect 26835 20349 26847 20352
rect 26789 20343 26847 20349
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 27065 20383 27123 20389
rect 27065 20349 27077 20383
rect 27111 20380 27123 20383
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 27111 20352 27261 20380
rect 27111 20349 27123 20352
rect 27065 20343 27123 20349
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 27341 20383 27399 20389
rect 27341 20349 27353 20383
rect 27387 20349 27399 20383
rect 27341 20343 27399 20349
rect 14599 20284 14780 20312
rect 27356 20312 27384 20343
rect 27430 20340 27436 20392
rect 27488 20340 27494 20392
rect 28994 20340 29000 20392
rect 29052 20340 29058 20392
rect 29089 20383 29147 20389
rect 29089 20349 29101 20383
rect 29135 20380 29147 20383
rect 29273 20383 29331 20389
rect 29273 20380 29285 20383
rect 29135 20352 29285 20380
rect 29135 20349 29147 20352
rect 29089 20343 29147 20349
rect 29273 20349 29285 20352
rect 29319 20349 29331 20383
rect 29273 20343 29331 20349
rect 29365 20383 29423 20389
rect 29365 20349 29377 20383
rect 29411 20380 29423 20383
rect 29549 20383 29607 20389
rect 29549 20380 29561 20383
rect 29411 20352 29561 20380
rect 29411 20349 29423 20352
rect 29365 20343 29423 20349
rect 29549 20349 29561 20352
rect 29595 20349 29607 20383
rect 29549 20343 29607 20349
rect 27525 20315 27583 20321
rect 27525 20312 27537 20315
rect 27356 20284 27537 20312
rect 14599 20281 14611 20284
rect 14553 20275 14611 20281
rect 27525 20281 27537 20284
rect 27571 20281 27583 20315
rect 27525 20275 27583 20281
rect 11747 20216 12572 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14332 20216 14841 20244
rect 14332 20204 14338 20216
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 14829 20207 14887 20213
rect 16114 20204 16120 20256
rect 16172 20204 16178 20256
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 19058 20244 19064 20256
rect 18831 20216 19064 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 21450 20204 21456 20256
rect 21508 20204 21514 20256
rect 26694 20204 26700 20256
rect 26752 20204 26758 20256
rect 552 20154 31648 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 12096 20154
rect 12148 20102 12160 20154
rect 12212 20102 12224 20154
rect 12276 20102 12288 20154
rect 12340 20102 12352 20154
rect 12404 20102 19870 20154
rect 19922 20102 19934 20154
rect 19986 20102 19998 20154
rect 20050 20102 20062 20154
rect 20114 20102 20126 20154
rect 20178 20102 27644 20154
rect 27696 20102 27708 20154
rect 27760 20102 27772 20154
rect 27824 20102 27836 20154
rect 27888 20102 27900 20154
rect 27952 20102 31648 20154
rect 552 20080 31648 20102
rect 1118 20000 1124 20052
rect 1176 20000 1182 20052
rect 1394 20000 1400 20052
rect 1452 20000 1458 20052
rect 3326 20000 3332 20052
rect 3384 20000 3390 20052
rect 6454 20000 6460 20052
rect 6512 20000 6518 20052
rect 11238 20000 11244 20052
rect 11296 20040 11302 20052
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 11296 20012 11713 20040
rect 11296 20000 11302 20012
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 17310 20000 17316 20052
rect 17368 20040 17374 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 17368 20012 17693 20040
rect 17368 20000 17374 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 19702 20000 19708 20052
rect 19760 20000 19766 20052
rect 24213 20043 24271 20049
rect 24213 20009 24225 20043
rect 24259 20040 24271 20043
rect 24394 20040 24400 20052
rect 24259 20012 24400 20040
rect 24259 20009 24271 20012
rect 24213 20003 24271 20009
rect 24394 20000 24400 20012
rect 24452 20000 24458 20052
rect 2501 19975 2559 19981
rect 2501 19941 2513 19975
rect 2547 19972 2559 19975
rect 3605 19975 3663 19981
rect 2547 19944 2728 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 1210 19864 1216 19916
rect 1268 19864 1274 19916
rect 1486 19864 1492 19916
rect 1544 19864 1550 19916
rect 1762 19864 1768 19916
rect 1820 19864 1826 19916
rect 2700 19913 2728 19944
rect 3605 19941 3617 19975
rect 3651 19972 3663 19975
rect 4157 19975 4215 19981
rect 3651 19944 3832 19972
rect 3651 19941 3663 19944
rect 3605 19935 3663 19941
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 1949 19907 2007 19913
rect 1949 19873 1961 19907
rect 1995 19904 2007 19907
rect 2133 19907 2191 19913
rect 2133 19904 2145 19907
rect 1995 19876 2145 19904
rect 1995 19873 2007 19876
rect 1949 19867 2007 19873
rect 2133 19873 2145 19876
rect 2179 19873 2191 19907
rect 2133 19867 2191 19873
rect 2593 19907 2651 19913
rect 2593 19873 2605 19907
rect 2639 19873 2651 19907
rect 2593 19867 2651 19873
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 2961 19907 3019 19913
rect 2961 19904 2973 19907
rect 2823 19876 2973 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 2961 19873 2973 19876
rect 3007 19873 3019 19907
rect 2961 19867 3019 19873
rect 3053 19907 3111 19913
rect 3053 19873 3065 19907
rect 3099 19904 3111 19907
rect 3237 19907 3295 19913
rect 3237 19904 3249 19907
rect 3099 19876 3249 19904
rect 3099 19873 3111 19876
rect 3053 19867 3111 19873
rect 3237 19873 3249 19876
rect 3283 19873 3295 19907
rect 3237 19867 3295 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1872 19836 1900 19867
rect 1719 19808 1900 19836
rect 2608 19836 2636 19867
rect 3694 19864 3700 19916
rect 3752 19864 3758 19916
rect 3804 19913 3832 19944
rect 4157 19941 4169 19975
rect 4203 19972 4215 19975
rect 5261 19975 5319 19981
rect 4203 19944 4384 19972
rect 4203 19941 4215 19944
rect 4157 19935 4215 19941
rect 3789 19907 3847 19913
rect 3789 19873 3801 19907
rect 3835 19873 3847 19907
rect 3789 19867 3847 19873
rect 4246 19864 4252 19916
rect 4304 19864 4310 19916
rect 4356 19913 4384 19944
rect 5261 19941 5273 19975
rect 5307 19972 5319 19975
rect 6733 19975 6791 19981
rect 6733 19972 6745 19975
rect 5307 19944 5488 19972
rect 5307 19941 5319 19944
rect 5261 19935 5319 19941
rect 5460 19913 5488 19944
rect 6564 19944 6745 19972
rect 6564 19913 6592 19944
rect 6733 19941 6745 19944
rect 6779 19941 6791 19975
rect 8849 19975 8907 19981
rect 8849 19972 8861 19975
rect 6733 19935 6791 19941
rect 8680 19944 8861 19972
rect 8680 19913 8708 19944
rect 8849 19941 8861 19944
rect 8895 19941 8907 19975
rect 11425 19975 11483 19981
rect 11425 19972 11437 19975
rect 8849 19935 8907 19941
rect 11256 19944 11437 19972
rect 4341 19907 4399 19913
rect 4341 19873 4353 19907
rect 4387 19873 4399 19907
rect 4341 19867 4399 19873
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 4479 19876 4629 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4617 19873 4629 19876
rect 4663 19873 4675 19907
rect 4617 19867 4675 19873
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 4893 19907 4951 19913
rect 4893 19904 4905 19907
rect 4755 19876 4905 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 4893 19873 4905 19876
rect 4939 19873 4951 19907
rect 4893 19867 4951 19873
rect 5353 19907 5411 19913
rect 5353 19873 5365 19907
rect 5399 19873 5411 19907
rect 5353 19867 5411 19873
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5583 19876 6009 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 6549 19907 6607 19913
rect 6549 19873 6561 19907
rect 6595 19873 6607 19907
rect 6549 19867 6607 19873
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19873 6699 19907
rect 6641 19867 6699 19873
rect 8113 19907 8171 19913
rect 8113 19873 8125 19907
rect 8159 19904 8171 19907
rect 8297 19907 8355 19913
rect 8297 19904 8309 19907
rect 8159 19876 8309 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 8297 19873 8309 19876
rect 8343 19873 8355 19907
rect 8297 19867 8355 19873
rect 8389 19907 8447 19913
rect 8389 19873 8401 19907
rect 8435 19904 8447 19907
rect 8573 19907 8631 19913
rect 8573 19904 8585 19907
rect 8435 19876 8585 19904
rect 8435 19873 8447 19876
rect 8389 19867 8447 19873
rect 8573 19873 8585 19876
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 8665 19907 8723 19913
rect 8665 19873 8677 19907
rect 8711 19873 8723 19907
rect 8665 19867 8723 19873
rect 2866 19836 2872 19848
rect 2608 19808 2872 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 5368 19768 5396 19867
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19836 6147 19839
rect 6656 19836 6684 19867
rect 8754 19864 8760 19916
rect 8812 19864 8818 19916
rect 9582 19864 9588 19916
rect 9640 19864 9646 19916
rect 10318 19864 10324 19916
rect 10376 19864 10382 19916
rect 10594 19864 10600 19916
rect 10652 19864 10658 19916
rect 11256 19913 11284 19944
rect 11425 19941 11437 19944
rect 11471 19941 11483 19975
rect 11977 19975 12035 19981
rect 11977 19972 11989 19975
rect 11425 19935 11483 19941
rect 11808 19944 11989 19972
rect 11808 19913 11836 19944
rect 11977 19941 11989 19944
rect 12023 19941 12035 19975
rect 11977 19935 12035 19941
rect 13909 19975 13967 19981
rect 13909 19941 13921 19975
rect 13955 19972 13967 19975
rect 19153 19975 19211 19981
rect 19153 19972 19165 19975
rect 13955 19944 14412 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19873 11851 19907
rect 11793 19867 11851 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 6135 19808 6684 19836
rect 10689 19839 10747 19845
rect 6135 19805 6147 19808
rect 6089 19799 6147 19805
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 11348 19836 11376 19867
rect 10735 19808 11376 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 5534 19768 5540 19780
rect 5368 19740 5540 19768
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 11149 19771 11207 19777
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11900 19768 11928 19867
rect 12710 19864 12716 19916
rect 12768 19864 12774 19916
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 13219 19876 13369 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 13357 19873 13369 19876
rect 13403 19873 13415 19907
rect 13357 19867 13415 19873
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13633 19907 13691 19913
rect 13633 19904 13645 19907
rect 13495 19876 13645 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13633 19873 13645 19876
rect 13679 19873 13691 19907
rect 13633 19867 13691 19873
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 14001 19907 14059 19913
rect 14001 19873 14013 19907
rect 14047 19904 14059 19907
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 14047 19876 14197 19904
rect 14047 19873 14059 19876
rect 14001 19867 14059 19873
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 13740 19836 13768 19867
rect 14274 19864 14280 19916
rect 14332 19864 14338 19916
rect 14384 19913 14412 19944
rect 18984 19944 19165 19972
rect 14369 19907 14427 19913
rect 14369 19873 14381 19907
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15335 19876 15485 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15611 19876 15761 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 15841 19907 15899 19913
rect 15841 19873 15853 19907
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 13740 19808 14473 19836
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 15856 19836 15884 19867
rect 16114 19864 16120 19916
rect 16172 19864 16178 19916
rect 17218 19864 17224 19916
rect 17276 19864 17282 19916
rect 18984 19913 19012 19944
rect 19153 19941 19165 19944
rect 19199 19941 19211 19975
rect 20533 19975 20591 19981
rect 20533 19972 20545 19975
rect 19153 19935 19211 19941
rect 20088 19944 20545 19972
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19904 17463 19907
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 17451 19876 17601 19904
rect 17451 19873 17463 19876
rect 17405 19867 17463 19873
rect 17589 19873 17601 19876
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 18693 19907 18751 19913
rect 18693 19873 18705 19907
rect 18739 19904 18751 19907
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18739 19876 18889 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 15856 19808 16221 19836
rect 14461 19799 14519 19805
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17328 19836 17356 19867
rect 19058 19864 19064 19916
rect 19116 19864 19122 19916
rect 20088 19913 20116 19944
rect 20533 19941 20545 19944
rect 20579 19941 20591 19975
rect 26145 19975 26203 19981
rect 26145 19972 26157 19975
rect 20533 19935 20591 19941
rect 25976 19944 26157 19972
rect 19797 19907 19855 19913
rect 19797 19873 19809 19907
rect 19843 19904 19855 19907
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19843 19876 19993 19904
rect 19843 19873 19855 19876
rect 19797 19867 19855 19873
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20073 19907 20131 19913
rect 20073 19873 20085 19907
rect 20119 19873 20131 19907
rect 20073 19867 20131 19873
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20257 19907 20315 19913
rect 20257 19873 20269 19907
rect 20303 19904 20315 19907
rect 20441 19907 20499 19913
rect 20441 19904 20453 19907
rect 20303 19876 20453 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20441 19873 20453 19876
rect 20487 19873 20499 19907
rect 20441 19867 20499 19873
rect 21450 19864 21456 19916
rect 21508 19864 21514 19916
rect 25976 19913 26004 19944
rect 26145 19941 26157 19944
rect 26191 19941 26203 19975
rect 26145 19935 26203 19941
rect 28261 19975 28319 19981
rect 28261 19941 28273 19975
rect 28307 19972 28319 19975
rect 28307 19944 28488 19972
rect 28307 19941 28319 19944
rect 28261 19935 28319 19941
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19904 21603 19907
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21591 19876 21741 19904
rect 21591 19873 21603 19876
rect 21545 19867 21603 19873
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 21821 19907 21879 19913
rect 21821 19873 21833 19907
rect 21867 19904 21879 19907
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 21867 19876 22017 19904
rect 21867 19873 21879 19876
rect 21821 19867 21879 19873
rect 22005 19873 22017 19876
rect 22051 19873 22063 19907
rect 22005 19867 22063 19873
rect 22097 19907 22155 19913
rect 22097 19873 22109 19907
rect 22143 19904 22155 19907
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 22143 19876 22293 19904
rect 22143 19873 22155 19876
rect 22097 19867 22155 19873
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22373 19907 22431 19913
rect 22373 19873 22385 19907
rect 22419 19904 22431 19907
rect 22557 19907 22615 19913
rect 22557 19904 22569 19907
rect 22419 19876 22569 19904
rect 22419 19873 22431 19876
rect 22373 19867 22431 19873
rect 22557 19873 22569 19876
rect 22603 19873 22615 19907
rect 22557 19867 22615 19873
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19904 22707 19907
rect 22833 19907 22891 19913
rect 22833 19904 22845 19907
rect 22695 19876 22845 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 22833 19873 22845 19876
rect 22879 19873 22891 19907
rect 22833 19867 22891 19873
rect 22925 19907 22983 19913
rect 22925 19873 22937 19907
rect 22971 19904 22983 19907
rect 23109 19907 23167 19913
rect 23109 19904 23121 19907
rect 22971 19876 23121 19904
rect 22971 19873 22983 19876
rect 22925 19867 22983 19873
rect 23109 19873 23121 19876
rect 23155 19873 23167 19907
rect 23109 19867 23167 19873
rect 24305 19907 24363 19913
rect 24305 19873 24317 19907
rect 24351 19904 24363 19907
rect 24489 19907 24547 19913
rect 24489 19904 24501 19907
rect 24351 19876 24501 19904
rect 24351 19873 24363 19876
rect 24305 19867 24363 19873
rect 24489 19873 24501 19876
rect 24535 19873 24547 19907
rect 24489 19867 24547 19873
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24765 19907 24823 19913
rect 24765 19904 24777 19907
rect 24627 19876 24777 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24765 19873 24777 19876
rect 24811 19873 24823 19907
rect 24765 19867 24823 19873
rect 24857 19907 24915 19913
rect 24857 19873 24869 19907
rect 24903 19904 24915 19907
rect 25041 19907 25099 19913
rect 25041 19904 25053 19907
rect 24903 19876 25053 19904
rect 24903 19873 24915 19876
rect 24857 19867 24915 19873
rect 25041 19873 25053 19876
rect 25087 19873 25099 19907
rect 25041 19867 25099 19873
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19904 25191 19907
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 25179 19876 25329 19904
rect 25179 19873 25191 19876
rect 25133 19867 25191 19873
rect 25317 19873 25329 19876
rect 25363 19873 25375 19907
rect 25317 19867 25375 19873
rect 25409 19907 25467 19913
rect 25409 19873 25421 19907
rect 25455 19904 25467 19907
rect 25593 19907 25651 19913
rect 25593 19904 25605 19907
rect 25455 19876 25605 19904
rect 25455 19873 25467 19876
rect 25409 19867 25467 19873
rect 25593 19873 25605 19876
rect 25639 19873 25651 19907
rect 25593 19867 25651 19873
rect 25685 19907 25743 19913
rect 25685 19873 25697 19907
rect 25731 19904 25743 19907
rect 25869 19907 25927 19913
rect 25869 19904 25881 19907
rect 25731 19876 25881 19904
rect 25731 19873 25743 19876
rect 25685 19867 25743 19873
rect 25869 19873 25881 19876
rect 25915 19873 25927 19907
rect 25869 19867 25927 19873
rect 25961 19907 26019 19913
rect 25961 19873 25973 19907
rect 26007 19873 26019 19907
rect 25961 19867 26019 19873
rect 26050 19864 26056 19916
rect 26108 19864 26114 19916
rect 26605 19907 26663 19913
rect 26605 19873 26617 19907
rect 26651 19904 26663 19907
rect 26789 19907 26847 19913
rect 26789 19904 26801 19907
rect 26651 19876 26801 19904
rect 26651 19873 26663 19876
rect 26605 19867 26663 19873
rect 26789 19873 26801 19876
rect 26835 19873 26847 19907
rect 26789 19867 26847 19873
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19904 26939 19907
rect 27065 19907 27123 19913
rect 27065 19904 27077 19907
rect 26927 19876 27077 19904
rect 26927 19873 26939 19876
rect 26881 19867 26939 19873
rect 27065 19873 27077 19876
rect 27111 19873 27123 19907
rect 27065 19867 27123 19873
rect 27157 19907 27215 19913
rect 27157 19873 27169 19907
rect 27203 19873 27215 19907
rect 27157 19867 27215 19873
rect 17175 19808 17356 19836
rect 27172 19836 27200 19867
rect 27246 19864 27252 19916
rect 27304 19864 27310 19916
rect 28350 19864 28356 19916
rect 28408 19864 28414 19916
rect 28460 19913 28488 19944
rect 28445 19907 28503 19913
rect 28445 19873 28457 19907
rect 28491 19873 28503 19907
rect 28445 19867 28503 19873
rect 28537 19907 28595 19913
rect 28537 19873 28549 19907
rect 28583 19904 28595 19907
rect 28721 19907 28779 19913
rect 28721 19904 28733 19907
rect 28583 19876 28733 19904
rect 28583 19873 28595 19876
rect 28537 19867 28595 19873
rect 28721 19873 28733 19876
rect 28767 19873 28779 19907
rect 28721 19867 28779 19873
rect 28813 19907 28871 19913
rect 28813 19873 28825 19907
rect 28859 19904 28871 19907
rect 28997 19907 29055 19913
rect 28997 19904 29009 19907
rect 28859 19876 29009 19904
rect 28859 19873 28871 19876
rect 28813 19867 28871 19873
rect 28997 19873 29009 19876
rect 29043 19873 29055 19907
rect 28997 19867 29055 19873
rect 29089 19907 29147 19913
rect 29089 19873 29101 19907
rect 29135 19904 29147 19907
rect 29273 19907 29331 19913
rect 29273 19904 29285 19907
rect 29135 19876 29285 19904
rect 29135 19873 29147 19876
rect 29089 19867 29147 19873
rect 29273 19873 29285 19876
rect 29319 19873 29331 19907
rect 29273 19867 29331 19873
rect 29365 19907 29423 19913
rect 29365 19873 29377 19907
rect 29411 19904 29423 19907
rect 29549 19907 29607 19913
rect 29549 19904 29561 19907
rect 29411 19876 29561 19904
rect 29411 19873 29423 19876
rect 29365 19867 29423 19873
rect 29549 19873 29561 19876
rect 29595 19873 29607 19907
rect 29549 19867 29607 19873
rect 27341 19839 27399 19845
rect 27341 19836 27353 19839
rect 27172 19808 27353 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 27341 19805 27353 19808
rect 27387 19805 27399 19839
rect 27341 19799 27399 19805
rect 11195 19740 11928 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 2225 19703 2283 19709
rect 2225 19669 2237 19703
rect 2271 19700 2283 19703
rect 2774 19700 2780 19712
rect 2271 19672 2780 19700
rect 2271 19669 2283 19672
rect 2225 19663 2283 19669
rect 2774 19660 2780 19672
rect 2832 19660 2838 19712
rect 3881 19703 3939 19709
rect 3881 19669 3893 19703
rect 3927 19700 3939 19703
rect 4338 19700 4344 19712
rect 3927 19672 4344 19700
rect 3927 19669 3939 19672
rect 3881 19663 3939 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 4985 19703 5043 19709
rect 4985 19669 4997 19703
rect 5031 19700 5043 19703
rect 5442 19700 5448 19712
rect 5031 19672 5448 19700
rect 5031 19669 5043 19672
rect 4985 19663 5043 19669
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8386 19700 8392 19712
rect 8067 19672 8392 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 9677 19703 9735 19709
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 9766 19700 9772 19712
rect 9723 19672 9772 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10413 19703 10471 19709
rect 10413 19669 10425 19703
rect 10459 19700 10471 19703
rect 10502 19700 10508 19712
rect 10459 19672 10508 19700
rect 10459 19669 10471 19672
rect 10413 19663 10471 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 12618 19660 12624 19712
rect 12676 19660 12682 19712
rect 12986 19660 12992 19712
rect 13044 19700 13050 19712
rect 13081 19703 13139 19709
rect 13081 19700 13093 19703
rect 13044 19672 13093 19700
rect 13044 19660 13050 19672
rect 13081 19669 13093 19672
rect 13127 19669 13139 19703
rect 13081 19663 13139 19669
rect 15194 19660 15200 19712
rect 15252 19660 15258 19712
rect 18598 19660 18604 19712
rect 18656 19660 18662 19712
rect 22830 19660 22836 19712
rect 22888 19700 22894 19712
rect 23201 19703 23259 19709
rect 23201 19700 23213 19703
rect 22888 19672 23213 19700
rect 22888 19660 22894 19672
rect 23201 19669 23213 19672
rect 23247 19669 23259 19703
rect 23201 19663 23259 19669
rect 26510 19660 26516 19712
rect 26568 19660 26574 19712
rect 29178 19660 29184 19712
rect 29236 19700 29242 19712
rect 29641 19703 29699 19709
rect 29641 19700 29653 19703
rect 29236 19672 29653 19700
rect 29236 19660 29242 19672
rect 29641 19669 29653 19672
rect 29687 19669 29699 19703
rect 29641 19663 29699 19669
rect 552 19610 31648 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 11436 19610
rect 11488 19558 11500 19610
rect 11552 19558 11564 19610
rect 11616 19558 11628 19610
rect 11680 19558 11692 19610
rect 11744 19558 19210 19610
rect 19262 19558 19274 19610
rect 19326 19558 19338 19610
rect 19390 19558 19402 19610
rect 19454 19558 19466 19610
rect 19518 19558 26984 19610
rect 27036 19558 27048 19610
rect 27100 19558 27112 19610
rect 27164 19558 27176 19610
rect 27228 19558 27240 19610
rect 27292 19558 31648 19610
rect 552 19536 31648 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2133 19499 2191 19505
rect 2133 19496 2145 19499
rect 1544 19468 2145 19496
rect 1544 19456 1550 19468
rect 2133 19465 2145 19468
rect 2179 19465 2191 19499
rect 2133 19459 2191 19465
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 4304 19468 4445 19496
rect 4304 19456 4310 19468
rect 4433 19465 4445 19468
rect 4479 19465 4491 19499
rect 4433 19459 4491 19465
rect 8849 19499 8907 19505
rect 8849 19465 8861 19499
rect 8895 19496 8907 19499
rect 9582 19496 9588 19508
rect 8895 19468 9588 19496
rect 8895 19465 8907 19468
rect 8849 19459 8907 19465
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 10137 19499 10195 19505
rect 10137 19465 10149 19499
rect 10183 19496 10195 19499
rect 10318 19496 10324 19508
rect 10183 19468 10324 19496
rect 10183 19465 10195 19468
rect 10137 19459 10195 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10594 19456 10600 19508
rect 10652 19456 10658 19508
rect 12710 19456 12716 19508
rect 12768 19496 12774 19508
rect 12805 19499 12863 19505
rect 12805 19496 12817 19499
rect 12768 19468 12817 19496
rect 12768 19456 12774 19468
rect 12805 19465 12817 19468
rect 12851 19465 12863 19499
rect 12805 19459 12863 19465
rect 17218 19456 17224 19508
rect 17276 19496 17282 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17276 19468 17877 19496
rect 17276 19456 17282 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 20162 19456 20168 19508
rect 20220 19456 20226 19508
rect 25593 19499 25651 19505
rect 25593 19465 25605 19499
rect 25639 19496 25651 19499
rect 26050 19496 26056 19508
rect 25639 19468 26056 19496
rect 25639 19465 25651 19468
rect 25593 19459 25651 19465
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 26605 19499 26663 19505
rect 26605 19465 26617 19499
rect 26651 19496 26663 19499
rect 27338 19496 27344 19508
rect 26651 19468 27344 19496
rect 26651 19465 26663 19468
rect 26605 19459 26663 19465
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 28350 19456 28356 19508
rect 28408 19496 28414 19508
rect 28721 19499 28779 19505
rect 28721 19496 28733 19499
rect 28408 19468 28733 19496
rect 28408 19456 28414 19468
rect 28721 19465 28733 19468
rect 28767 19465 28779 19499
rect 28721 19459 28779 19465
rect 28994 19456 29000 19508
rect 29052 19496 29058 19508
rect 29089 19499 29147 19505
rect 29089 19496 29101 19499
rect 29052 19468 29101 19496
rect 29052 19456 29058 19468
rect 29089 19465 29101 19468
rect 29135 19465 29147 19499
rect 29089 19459 29147 19465
rect 23017 19431 23075 19437
rect 23017 19397 23029 19431
rect 23063 19428 23075 19431
rect 23063 19400 23336 19428
rect 23063 19397 23075 19400
rect 23017 19391 23075 19397
rect 12618 19360 12624 19372
rect 12268 19332 12624 19360
rect 1486 19252 1492 19304
rect 1544 19252 1550 19304
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19292 1639 19295
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1627 19264 1777 19292
rect 1627 19261 1639 19264
rect 1581 19255 1639 19261
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 2041 19295 2099 19301
rect 2041 19292 2053 19295
rect 1903 19264 2053 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 2041 19261 2053 19264
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 2774 19252 2780 19304
rect 2832 19252 2838 19304
rect 2866 19252 2872 19304
rect 2924 19252 2930 19304
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 3697 19295 3755 19301
rect 3697 19292 3709 19295
rect 3568 19264 3709 19292
rect 3568 19252 3574 19264
rect 3697 19261 3709 19264
rect 3743 19261 3755 19295
rect 3697 19255 3755 19261
rect 4338 19252 4344 19304
rect 4396 19252 4402 19304
rect 5442 19252 5448 19304
rect 5500 19252 5506 19304
rect 5534 19252 5540 19304
rect 5592 19252 5598 19304
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7699 19264 7849 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 7837 19255 7895 19261
rect 7929 19295 7987 19301
rect 7929 19261 7941 19295
rect 7975 19292 7987 19295
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 7975 19264 8125 19292
rect 7975 19261 7987 19264
rect 7929 19255 7987 19261
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8113 19255 8171 19261
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 8220 19224 8248 19255
rect 8386 19252 8392 19304
rect 8444 19252 8450 19304
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 9125 19295 9183 19301
rect 9125 19292 9137 19295
rect 8987 19264 9137 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 9125 19261 9137 19264
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 8481 19227 8539 19233
rect 8481 19224 8493 19227
rect 8220 19196 8493 19224
rect 8481 19193 8493 19196
rect 8527 19193 8539 19227
rect 9232 19224 9260 19255
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 9907 19264 10057 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10045 19255 10103 19261
rect 10502 19252 10508 19304
rect 10560 19252 10566 19304
rect 12268 19301 12296 19332
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 15580 19332 15792 19360
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19261 12403 19295
rect 12345 19255 12403 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 9401 19227 9459 19233
rect 9401 19224 9413 19227
rect 9232 19196 9413 19224
rect 8481 19187 8539 19193
rect 9401 19193 9413 19196
rect 9447 19193 9459 19227
rect 9401 19187 9459 19193
rect 12161 19227 12219 19233
rect 12161 19193 12173 19227
rect 12207 19224 12219 19227
rect 12360 19224 12388 19255
rect 12207 19196 12388 19224
rect 12912 19224 12940 19255
rect 12986 19252 12992 19304
rect 13044 19252 13050 19304
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13127 19264 13553 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 13633 19227 13691 19233
rect 13633 19224 13645 19227
rect 12912 19196 13645 19224
rect 12207 19193 12219 19196
rect 12161 19187 12219 19193
rect 13633 19193 13645 19196
rect 13679 19193 13691 19227
rect 15028 19224 15056 19255
rect 15194 19252 15200 19304
rect 15252 19252 15258 19304
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15580 19292 15608 19332
rect 15764 19301 15792 19332
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18656 19332 19288 19360
rect 18656 19320 18662 19332
rect 15335 19264 15608 19292
rect 15657 19295 15715 19301
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19261 15807 19295
rect 15749 19255 15807 19261
rect 15565 19227 15623 19233
rect 15565 19224 15577 19227
rect 15028 19196 15577 19224
rect 13633 19187 13691 19193
rect 15565 19193 15577 19196
rect 15611 19193 15623 19227
rect 15672 19224 15700 19255
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 19260 19301 19288 19332
rect 23032 19332 23244 19360
rect 17221 19295 17279 19301
rect 17221 19261 17233 19295
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 17359 19264 17509 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 17773 19295 17831 19301
rect 17773 19292 17785 19295
rect 17635 19264 17785 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 17773 19261 17785 19264
rect 17819 19261 17831 19295
rect 17773 19255 17831 19261
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18923 19264 19073 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 19153 19295 19211 19301
rect 19153 19261 19165 19295
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 20257 19295 20315 19301
rect 20257 19261 20269 19295
rect 20303 19292 20315 19295
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 20303 19264 20453 19292
rect 20303 19261 20315 19264
rect 20257 19255 20315 19261
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 20579 19264 20668 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 15672 19196 15853 19224
rect 15565 19187 15623 19193
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15841 19187 15899 19193
rect 17037 19227 17095 19233
rect 17037 19193 17049 19227
rect 17083 19224 17095 19227
rect 17236 19224 17264 19255
rect 17083 19196 17264 19224
rect 19168 19224 19196 19255
rect 19337 19227 19395 19233
rect 19337 19224 19349 19227
rect 19168 19196 19349 19224
rect 17083 19193 17095 19196
rect 17037 19187 17095 19193
rect 19337 19193 19349 19196
rect 19383 19193 19395 19227
rect 19337 19187 19395 19193
rect 3694 19116 3700 19168
rect 3752 19156 3758 19168
rect 3789 19159 3847 19165
rect 3789 19156 3801 19159
rect 3752 19128 3801 19156
rect 3752 19116 3758 19128
rect 3789 19125 3801 19128
rect 3835 19125 3847 19159
rect 3789 19119 3847 19125
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7561 19159 7619 19165
rect 7561 19156 7573 19159
rect 7340 19128 7573 19156
rect 7340 19116 7346 19128
rect 7561 19125 7573 19128
rect 7607 19125 7619 19159
rect 7561 19119 7619 19125
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 14921 19159 14979 19165
rect 14921 19156 14933 19159
rect 14700 19128 14933 19156
rect 14700 19116 14706 19128
rect 14921 19125 14933 19128
rect 14967 19125 14979 19159
rect 14921 19119 14979 19125
rect 18782 19116 18788 19168
rect 18840 19116 18846 19168
rect 20640 19156 20668 19264
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 20717 19227 20775 19233
rect 20717 19193 20729 19227
rect 20763 19224 20775 19227
rect 20916 19224 20944 19255
rect 22830 19252 22836 19304
rect 22888 19252 22894 19304
rect 20763 19196 20944 19224
rect 22741 19227 22799 19233
rect 20763 19193 20775 19196
rect 20717 19187 20775 19193
rect 22741 19193 22753 19227
rect 22787 19224 22799 19227
rect 23032 19224 23060 19332
rect 23216 19301 23244 19332
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 23201 19295 23259 19301
rect 23201 19261 23213 19295
rect 23247 19261 23259 19295
rect 23308 19292 23336 19400
rect 23477 19295 23535 19301
rect 23477 19292 23489 19295
rect 23308 19264 23489 19292
rect 23201 19255 23259 19261
rect 23477 19261 23489 19264
rect 23523 19261 23535 19295
rect 23477 19255 23535 19261
rect 25685 19295 25743 19301
rect 25685 19261 25697 19295
rect 25731 19292 25743 19295
rect 26510 19292 26516 19304
rect 25731 19264 26516 19292
rect 25731 19261 25743 19264
rect 25685 19255 25743 19261
rect 22787 19196 23060 19224
rect 23124 19224 23152 19255
rect 26510 19252 26516 19264
rect 26568 19252 26574 19304
rect 26694 19252 26700 19304
rect 26752 19252 26758 19304
rect 27982 19252 27988 19304
rect 28040 19292 28046 19304
rect 28077 19295 28135 19301
rect 28077 19292 28089 19295
rect 28040 19264 28089 19292
rect 28040 19252 28046 19264
rect 28077 19261 28089 19264
rect 28123 19261 28135 19295
rect 28077 19255 28135 19261
rect 28169 19295 28227 19301
rect 28169 19261 28181 19295
rect 28215 19292 28227 19295
rect 28353 19295 28411 19301
rect 28353 19292 28365 19295
rect 28215 19264 28365 19292
rect 28215 19261 28227 19264
rect 28169 19255 28227 19261
rect 28353 19261 28365 19264
rect 28399 19261 28411 19295
rect 28353 19255 28411 19261
rect 28445 19295 28503 19301
rect 28445 19261 28457 19295
rect 28491 19292 28503 19295
rect 28629 19295 28687 19301
rect 28629 19292 28641 19295
rect 28491 19264 28641 19292
rect 28491 19261 28503 19264
rect 28445 19255 28503 19261
rect 28629 19261 28641 19264
rect 28675 19261 28687 19295
rect 28629 19255 28687 19261
rect 29178 19252 29184 19304
rect 29236 19252 29242 19304
rect 23293 19227 23351 19233
rect 23293 19224 23305 19227
rect 23124 19196 23305 19224
rect 22787 19193 22799 19196
rect 22741 19187 22799 19193
rect 23293 19193 23305 19196
rect 23339 19193 23351 19227
rect 23293 19187 23351 19193
rect 20993 19159 21051 19165
rect 20993 19156 21005 19159
rect 20640 19128 21005 19156
rect 20993 19125 21005 19128
rect 21039 19125 21051 19159
rect 20993 19119 21051 19125
rect 23382 19116 23388 19168
rect 23440 19156 23446 19168
rect 23569 19159 23627 19165
rect 23569 19156 23581 19159
rect 23440 19128 23581 19156
rect 23440 19116 23446 19128
rect 23569 19125 23581 19128
rect 23615 19125 23627 19159
rect 23569 19119 23627 19125
rect 552 19066 31648 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31648 19066
rect 552 18992 31648 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1544 18924 1593 18952
rect 1544 18912 1550 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 3510 18912 3516 18964
rect 3568 18912 3574 18964
rect 9217 18955 9275 18961
rect 9217 18921 9229 18955
rect 9263 18952 9275 18955
rect 9306 18952 9312 18964
rect 9263 18924 9312 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 17126 18912 17132 18964
rect 17184 18952 17190 18964
rect 17773 18955 17831 18961
rect 17773 18952 17785 18955
rect 17184 18924 17785 18952
rect 17184 18912 17190 18924
rect 17773 18921 17785 18924
rect 17819 18921 17831 18955
rect 17773 18915 17831 18921
rect 20806 18912 20812 18964
rect 20864 18912 20870 18964
rect 27982 18912 27988 18964
rect 28040 18912 28046 18964
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 1688 18856 2421 18884
rect 1688 18825 1716 18856
rect 2409 18853 2421 18856
rect 2455 18853 2467 18887
rect 6181 18887 6239 18893
rect 6181 18884 6193 18887
rect 2409 18847 2467 18853
rect 6012 18856 6193 18884
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 1762 18776 1768 18828
rect 1820 18776 1826 18828
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1903 18788 2053 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2317 18819 2375 18825
rect 2317 18816 2329 18819
rect 2179 18788 2329 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 2317 18785 2329 18788
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18816 3479 18819
rect 3510 18816 3516 18828
rect 3467 18788 3516 18816
rect 3467 18785 3479 18788
rect 3421 18779 3479 18785
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 3694 18776 3700 18828
rect 3752 18776 3758 18828
rect 6012 18825 6040 18856
rect 6181 18853 6193 18856
rect 6227 18853 6239 18887
rect 8297 18887 8355 18893
rect 8297 18884 8309 18887
rect 6181 18847 6239 18853
rect 8128 18856 8309 18884
rect 3789 18819 3847 18825
rect 3789 18785 3801 18819
rect 3835 18816 3847 18819
rect 3973 18819 4031 18825
rect 3973 18816 3985 18819
rect 3835 18788 3985 18816
rect 3835 18785 3847 18788
rect 3789 18779 3847 18785
rect 3973 18785 3985 18788
rect 4019 18785 4031 18819
rect 3973 18779 4031 18785
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4111 18788 4261 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18816 4399 18819
rect 4525 18819 4583 18825
rect 4525 18816 4537 18819
rect 4387 18788 4537 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4525 18785 4537 18788
rect 4571 18785 4583 18819
rect 4525 18779 4583 18785
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 4801 18819 4859 18825
rect 4801 18816 4813 18819
rect 4663 18788 4813 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 4801 18785 4813 18788
rect 4847 18785 4859 18819
rect 4801 18779 4859 18785
rect 4893 18819 4951 18825
rect 4893 18785 4905 18819
rect 4939 18816 4951 18819
rect 5077 18819 5135 18825
rect 5077 18816 5089 18819
rect 4939 18788 5089 18816
rect 4939 18785 4951 18788
rect 4893 18779 4951 18785
rect 5077 18785 5089 18788
rect 5123 18785 5135 18819
rect 5077 18779 5135 18785
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 5215 18788 5365 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5353 18785 5365 18788
rect 5399 18785 5411 18819
rect 5353 18779 5411 18785
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 6104 18748 6132 18779
rect 7282 18776 7288 18828
rect 7340 18776 7346 18828
rect 8128 18825 8156 18856
rect 8297 18853 8309 18856
rect 8343 18853 8355 18887
rect 8297 18847 8355 18853
rect 9861 18887 9919 18893
rect 9861 18853 9873 18887
rect 9907 18884 9919 18887
rect 12434 18884 12440 18896
rect 9907 18856 10088 18884
rect 9907 18853 9919 18856
rect 9861 18847 9919 18853
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7607 18788 7757 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7883 18788 8033 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 9309 18819 9367 18825
rect 9309 18785 9321 18819
rect 9355 18816 9367 18819
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 9355 18788 9505 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18785 9643 18819
rect 9585 18779 9643 18785
rect 5491 18720 6132 18748
rect 7193 18751 7251 18757
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 8220 18748 8248 18779
rect 7239 18720 8248 18748
rect 9600 18748 9628 18779
rect 9950 18776 9956 18828
rect 10008 18776 10014 18828
rect 10060 18825 10088 18856
rect 12268 18856 12440 18884
rect 12268 18825 12296 18856
rect 12434 18844 12440 18856
rect 12492 18844 12498 18896
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 13096 18856 13277 18884
rect 13096 18825 13124 18856
rect 13265 18853 13277 18856
rect 13311 18853 13323 18887
rect 13265 18847 13323 18853
rect 14553 18887 14611 18893
rect 14553 18853 14565 18887
rect 14599 18884 14611 18887
rect 19521 18887 19579 18893
rect 19521 18884 19533 18887
rect 14599 18856 15608 18884
rect 14599 18853 14611 18856
rect 14553 18847 14611 18853
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12805 18819 12863 18825
rect 12805 18785 12817 18819
rect 12851 18816 12863 18819
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12851 18788 13001 18816
rect 12851 18785 12863 18788
rect 12805 18779 12863 18785
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13081 18819 13139 18825
rect 13081 18785 13093 18819
rect 13127 18785 13139 18819
rect 13081 18779 13139 18785
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 9600 18720 10149 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18748 12219 18751
rect 12360 18748 12388 18779
rect 12207 18720 12388 18748
rect 12437 18751 12495 18757
rect 12207 18717 12219 18720
rect 12161 18711 12219 18717
rect 12437 18717 12449 18751
rect 12483 18748 12495 18751
rect 13188 18748 13216 18779
rect 14642 18776 14648 18828
rect 14700 18776 14706 18828
rect 15580 18825 15608 18856
rect 19352 18856 19533 18884
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18816 14979 18819
rect 15105 18819 15163 18825
rect 15105 18816 15117 18819
rect 14967 18788 15117 18816
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 15105 18785 15117 18788
rect 15151 18785 15163 18819
rect 15105 18779 15163 18785
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 15381 18819 15439 18825
rect 15381 18816 15393 18819
rect 15243 18788 15393 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 15381 18785 15393 18788
rect 15427 18785 15439 18819
rect 15381 18779 15439 18785
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18785 15531 18819
rect 15473 18779 15531 18785
rect 15565 18819 15623 18825
rect 15565 18785 15577 18819
rect 15611 18785 15623 18819
rect 15565 18779 15623 18785
rect 12483 18720 13216 18748
rect 15488 18748 15516 18779
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 16853 18819 16911 18825
rect 16853 18816 16865 18819
rect 16724 18788 16865 18816
rect 16724 18776 16730 18788
rect 16853 18785 16865 18788
rect 16899 18785 16911 18819
rect 16853 18779 16911 18785
rect 16945 18819 17003 18825
rect 16945 18785 16957 18819
rect 16991 18816 17003 18819
rect 17129 18819 17187 18825
rect 17129 18816 17141 18819
rect 16991 18788 17141 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 17129 18785 17141 18788
rect 17175 18785 17187 18819
rect 17129 18779 17187 18785
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 17267 18788 17417 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17543 18788 17693 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 18782 18776 18788 18828
rect 18840 18776 18846 18828
rect 19352 18825 19380 18856
rect 19521 18853 19533 18856
rect 19567 18853 19579 18887
rect 21361 18887 21419 18893
rect 21361 18884 21373 18887
rect 19521 18847 19579 18853
rect 20916 18856 21373 18884
rect 20916 18825 20944 18856
rect 21361 18853 21373 18856
rect 21407 18853 21419 18887
rect 21361 18847 21419 18853
rect 23293 18887 23351 18893
rect 23293 18853 23305 18887
rect 23339 18884 23351 18887
rect 23339 18856 23520 18884
rect 23339 18853 23351 18856
rect 23293 18847 23351 18853
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18816 19119 18819
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 19107 18788 19257 18816
rect 19107 18785 19119 18788
rect 19061 18779 19119 18785
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 19429 18819 19487 18825
rect 19429 18785 19441 18819
rect 19475 18785 19487 18819
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 19429 18779 19487 18785
rect 20456 18788 20637 18816
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15488 18720 15669 18748
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 19444 18748 19472 18779
rect 18739 18720 19472 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 20456 18680 20484 18788
rect 20625 18785 20637 18788
rect 20671 18785 20683 18819
rect 20625 18779 20683 18785
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 21269 18819 21327 18825
rect 21269 18785 21281 18819
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18748 20591 18751
rect 21284 18748 21312 18779
rect 21542 18776 21548 18828
rect 21600 18776 21606 18828
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 21821 18819 21879 18825
rect 21821 18816 21833 18819
rect 21683 18788 21833 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 21821 18785 21833 18788
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 23382 18776 23388 18828
rect 23440 18776 23446 18828
rect 23492 18825 23520 18856
rect 23477 18819 23535 18825
rect 23477 18785 23489 18819
rect 23523 18785 23535 18819
rect 23477 18779 23535 18785
rect 23569 18819 23627 18825
rect 23569 18785 23581 18819
rect 23615 18816 23627 18819
rect 23753 18819 23811 18825
rect 23753 18816 23765 18819
rect 23615 18788 23765 18816
rect 23615 18785 23627 18788
rect 23569 18779 23627 18785
rect 23753 18785 23765 18788
rect 23799 18785 23811 18819
rect 23753 18779 23811 18785
rect 23845 18819 23903 18825
rect 23845 18785 23857 18819
rect 23891 18816 23903 18819
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23891 18788 24041 18816
rect 23891 18785 23903 18788
rect 23845 18779 23903 18785
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24029 18779 24087 18785
rect 24121 18819 24179 18825
rect 24121 18785 24133 18819
rect 24167 18816 24179 18819
rect 24305 18819 24363 18825
rect 24305 18816 24317 18819
rect 24167 18788 24317 18816
rect 24167 18785 24179 18788
rect 24121 18779 24179 18785
rect 24305 18785 24317 18788
rect 24351 18785 24363 18819
rect 24305 18779 24363 18785
rect 24397 18819 24455 18825
rect 24397 18785 24409 18819
rect 24443 18816 24455 18819
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24443 18788 24593 18816
rect 24443 18785 24455 18788
rect 24397 18779 24455 18785
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 24673 18819 24731 18825
rect 24673 18785 24685 18819
rect 24719 18816 24731 18819
rect 24857 18819 24915 18825
rect 24857 18816 24869 18819
rect 24719 18788 24869 18816
rect 24719 18785 24731 18788
rect 24673 18779 24731 18785
rect 24857 18785 24869 18788
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 24949 18819 25007 18825
rect 24949 18785 24961 18819
rect 24995 18816 25007 18819
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 24995 18788 25145 18816
rect 24995 18785 25007 18788
rect 24949 18779 25007 18785
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25409 18819 25467 18825
rect 25409 18816 25421 18819
rect 25271 18788 25421 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 25409 18785 25421 18788
rect 25455 18785 25467 18819
rect 25409 18779 25467 18785
rect 25501 18819 25559 18825
rect 25501 18785 25513 18819
rect 25547 18816 25559 18819
rect 25685 18819 25743 18825
rect 25685 18816 25697 18819
rect 25547 18788 25697 18816
rect 25547 18785 25559 18788
rect 25501 18779 25559 18785
rect 25685 18785 25697 18788
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 28077 18819 28135 18825
rect 28077 18785 28089 18819
rect 28123 18816 28135 18819
rect 28261 18819 28319 18825
rect 28261 18816 28273 18819
rect 28123 18788 28273 18816
rect 28123 18785 28135 18788
rect 28077 18779 28135 18785
rect 28261 18785 28273 18788
rect 28307 18785 28319 18819
rect 28261 18779 28319 18785
rect 28353 18819 28411 18825
rect 28353 18785 28365 18819
rect 28399 18785 28411 18819
rect 28353 18779 28411 18785
rect 20579 18720 21312 18748
rect 28368 18748 28396 18779
rect 28442 18776 28448 18828
rect 28500 18776 28506 18828
rect 28718 18776 28724 18828
rect 28776 18776 28782 18828
rect 28537 18751 28595 18757
rect 28537 18748 28549 18751
rect 28368 18720 28549 18748
rect 20579 18717 20591 18720
rect 20533 18711 20591 18717
rect 28537 18717 28549 18720
rect 28583 18717 28595 18751
rect 28537 18711 28595 18717
rect 21913 18683 21971 18689
rect 21913 18680 21925 18683
rect 20456 18652 21925 18680
rect 21913 18649 21925 18652
rect 21959 18649 21971 18683
rect 21913 18643 21971 18649
rect 5905 18615 5963 18621
rect 5905 18581 5917 18615
rect 5951 18612 5963 18615
rect 6546 18612 6552 18624
rect 5951 18584 6552 18612
rect 5951 18581 5963 18584
rect 5905 18575 5963 18581
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 7469 18615 7527 18621
rect 7469 18581 7481 18615
rect 7515 18612 7527 18615
rect 8018 18612 8024 18624
rect 7515 18584 8024 18612
rect 7515 18581 7527 18584
rect 7469 18575 7527 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14829 18615 14887 18621
rect 14829 18612 14841 18615
rect 14792 18584 14841 18612
rect 14792 18572 14798 18584
rect 14829 18581 14841 18584
rect 14875 18581 14887 18615
rect 14829 18575 14887 18581
rect 18874 18572 18880 18624
rect 18932 18612 18938 18624
rect 18969 18615 19027 18621
rect 18969 18612 18981 18615
rect 18932 18584 18981 18612
rect 18932 18572 18938 18584
rect 18969 18581 18981 18584
rect 19015 18581 19027 18615
rect 18969 18575 19027 18581
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 25777 18615 25835 18621
rect 25777 18612 25789 18615
rect 25648 18584 25789 18612
rect 25648 18572 25654 18584
rect 25777 18581 25789 18584
rect 25823 18581 25835 18615
rect 25777 18575 25835 18581
rect 28534 18572 28540 18624
rect 28592 18612 28598 18624
rect 28813 18615 28871 18621
rect 28813 18612 28825 18615
rect 28592 18584 28825 18612
rect 28592 18572 28598 18584
rect 28813 18581 28825 18584
rect 28859 18581 28871 18615
rect 28813 18575 28871 18581
rect 552 18522 31648 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31648 18522
rect 552 18448 31648 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 1762 18408 1768 18420
rect 1627 18380 1768 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 10008 18380 10701 18408
rect 10008 18368 10014 18380
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 10689 18371 10747 18377
rect 16666 18368 16672 18420
rect 16724 18368 16730 18420
rect 21177 18411 21235 18417
rect 21177 18377 21189 18411
rect 21223 18408 21235 18411
rect 21542 18408 21548 18420
rect 21223 18380 21548 18408
rect 21223 18377 21235 18380
rect 21177 18371 21235 18377
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 28353 18411 28411 18417
rect 28353 18377 28365 18411
rect 28399 18408 28411 18411
rect 28442 18408 28448 18420
rect 28399 18380 28448 18408
rect 28399 18377 28411 18380
rect 28353 18371 28411 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 28718 18368 28724 18420
rect 28776 18368 28782 18420
rect 10413 18343 10471 18349
rect 10413 18340 10425 18343
rect 9968 18312 10425 18340
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 3789 18275 3847 18281
rect 1903 18244 2084 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18173 1731 18207
rect 1673 18167 1731 18173
rect 1688 18136 1716 18167
rect 1946 18164 1952 18216
rect 2004 18164 2010 18216
rect 2056 18213 2084 18244
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 6641 18275 6699 18281
rect 6641 18272 6653 18275
rect 3835 18244 4016 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2317 18207 2375 18213
rect 2317 18204 2329 18207
rect 2179 18176 2329 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2317 18173 2329 18176
rect 2363 18173 2375 18207
rect 2317 18167 2375 18173
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2593 18207 2651 18213
rect 2593 18204 2605 18207
rect 2455 18176 2605 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2593 18173 2605 18176
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 2685 18139 2743 18145
rect 2685 18136 2697 18139
rect 1688 18108 2697 18136
rect 2685 18105 2697 18108
rect 2731 18105 2743 18139
rect 3620 18136 3648 18167
rect 3878 18164 3884 18216
rect 3936 18164 3942 18216
rect 3988 18213 4016 18244
rect 6472 18244 6653 18272
rect 6472 18213 6500 18244
rect 6641 18241 6653 18244
rect 6687 18241 6699 18275
rect 8113 18275 8171 18281
rect 8113 18272 8125 18275
rect 6641 18235 6699 18241
rect 7944 18244 8125 18272
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18173 4031 18207
rect 3973 18167 4031 18173
rect 4065 18207 4123 18213
rect 4065 18173 4077 18207
rect 4111 18204 4123 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4111 18176 4261 18204
rect 4111 18173 4123 18176
rect 4065 18167 4123 18173
rect 4249 18173 4261 18176
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18204 5963 18207
rect 6089 18207 6147 18213
rect 6089 18204 6101 18207
rect 5951 18176 6101 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 6089 18173 6101 18176
rect 6135 18173 6147 18207
rect 6089 18167 6147 18173
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 6227 18176 6377 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18173 6515 18207
rect 6457 18167 6515 18173
rect 6546 18164 6552 18216
rect 6604 18164 6610 18216
rect 7944 18213 7972 18244
rect 8113 18241 8125 18244
rect 8159 18241 8171 18275
rect 8113 18235 8171 18241
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18272 9367 18275
rect 9355 18244 9536 18272
rect 9355 18241 9367 18244
rect 9309 18235 9367 18241
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18204 7711 18207
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7699 18176 7849 18204
rect 7699 18173 7711 18176
rect 7653 18167 7711 18173
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 8018 18164 8024 18216
rect 8076 18164 8082 18216
rect 9508 18213 9536 18244
rect 9968 18213 9996 18312
rect 10413 18309 10425 18312
rect 10459 18309 10471 18343
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 10413 18303 10471 18309
rect 17052 18312 17785 18340
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18272 10195 18275
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 10183 18244 10640 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 10612 18213 10640 18244
rect 13280 18244 13645 18272
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18173 10011 18207
rect 9953 18167 10011 18173
rect 10045 18207 10103 18213
rect 10045 18173 10057 18207
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18173 10379 18207
rect 10321 18167 10379 18173
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 4341 18139 4399 18145
rect 4341 18136 4353 18139
rect 3620 18108 4353 18136
rect 2685 18099 2743 18105
rect 4341 18105 4353 18108
rect 4387 18105 4399 18139
rect 9416 18136 9444 18167
rect 9674 18136 9680 18148
rect 9416 18108 9680 18136
rect 4341 18099 4399 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 9861 18139 9919 18145
rect 9861 18105 9873 18139
rect 9907 18136 9919 18139
rect 10060 18136 10088 18167
rect 9907 18108 10088 18136
rect 9907 18105 9919 18108
rect 9861 18099 9919 18105
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 5813 18071 5871 18077
rect 5813 18068 5825 18071
rect 5684 18040 5825 18068
rect 5684 18028 5690 18040
rect 5813 18037 5825 18040
rect 5859 18037 5871 18071
rect 5813 18031 5871 18037
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 7524 18040 7573 18068
rect 7524 18028 7530 18040
rect 7561 18037 7573 18040
rect 7607 18037 7619 18071
rect 7561 18031 7619 18037
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18068 9643 18071
rect 10336 18068 10364 18167
rect 12710 18164 12716 18216
rect 12768 18164 12774 18216
rect 13280 18213 13308 18244
rect 13633 18241 13645 18244
rect 13679 18241 13691 18275
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 13633 18235 13691 18241
rect 15304 18244 15485 18272
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 13035 18176 13185 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18136 12679 18139
rect 13556 18136 13584 18167
rect 14734 18164 14740 18216
rect 14792 18164 14798 18216
rect 15304 18213 15332 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 17052 18213 17080 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 21453 18343 21511 18349
rect 21453 18309 21465 18343
rect 21499 18340 21511 18343
rect 21499 18312 22232 18340
rect 21499 18309 21511 18312
rect 21453 18303 21511 18309
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 19889 18275 19947 18281
rect 19889 18272 19901 18275
rect 17267 18244 17448 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17420 18213 17448 18244
rect 19444 18244 19901 18272
rect 15013 18207 15071 18213
rect 15013 18173 15025 18207
rect 15059 18204 15071 18207
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15059 18176 15209 18204
rect 15059 18173 15071 18176
rect 15013 18167 15071 18173
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15289 18167 15347 18173
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18204 16819 18207
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16807 18176 16957 18204
rect 16807 18173 16819 18176
rect 16761 18167 16819 18173
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18204 17555 18207
rect 17681 18207 17739 18213
rect 17681 18204 17693 18207
rect 17543 18176 17693 18204
rect 17543 18173 17555 18176
rect 17497 18167 17555 18173
rect 17681 18173 17693 18176
rect 17727 18173 17739 18207
rect 17681 18167 17739 18173
rect 12667 18108 13584 18136
rect 14645 18139 14703 18145
rect 12667 18105 12679 18108
rect 12621 18099 12679 18105
rect 14645 18105 14657 18139
rect 14691 18136 14703 18139
rect 15396 18136 15424 18167
rect 14691 18108 15424 18136
rect 14691 18105 14703 18108
rect 14645 18099 14703 18105
rect 9631 18040 10364 18068
rect 12897 18071 12955 18077
rect 9631 18037 9643 18040
rect 9585 18031 9643 18037
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13538 18068 13544 18080
rect 12943 18040 13544 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 14918 18028 14924 18080
rect 14976 18028 14982 18080
rect 17328 18068 17356 18167
rect 18874 18164 18880 18216
rect 18932 18164 18938 18216
rect 19444 18213 19472 18244
rect 19889 18241 19901 18244
rect 19935 18241 19947 18275
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 19889 18235 19947 18241
rect 21560 18244 22017 18272
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 19518 18164 19524 18216
rect 19576 18164 19582 18216
rect 21560 18213 21588 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 19613 18207 19671 18213
rect 19613 18173 19625 18207
rect 19659 18204 19671 18207
rect 19797 18207 19855 18213
rect 19797 18204 19809 18207
rect 19659 18176 19809 18204
rect 19659 18173 19671 18176
rect 19613 18167 19671 18173
rect 19797 18173 19809 18176
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 20073 18207 20131 18213
rect 20073 18173 20085 18207
rect 20119 18173 20131 18207
rect 20073 18167 20131 18173
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 21545 18207 21603 18213
rect 21545 18173 21557 18207
rect 21591 18173 21603 18207
rect 21545 18167 21603 18173
rect 19337 18139 19395 18145
rect 19337 18105 19349 18139
rect 19383 18136 19395 18139
rect 20088 18136 20116 18167
rect 19383 18108 20116 18136
rect 19383 18105 19395 18108
rect 19337 18099 19395 18105
rect 18046 18068 18052 18080
rect 17328 18040 18052 18068
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18966 18028 18972 18080
rect 19024 18028 19030 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 19668 18040 20177 18068
rect 19668 18028 19674 18040
rect 20165 18037 20177 18040
rect 20211 18037 20223 18071
rect 21284 18068 21312 18167
rect 21818 18164 21824 18216
rect 21876 18164 21882 18216
rect 22204 18213 22232 18312
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18272 25559 18275
rect 29917 18275 29975 18281
rect 29917 18272 29929 18275
rect 25547 18244 26096 18272
rect 25547 18241 25559 18244
rect 25501 18235 25559 18241
rect 21913 18207 21971 18213
rect 21913 18173 21925 18207
rect 21959 18173 21971 18207
rect 21913 18167 21971 18173
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18173 22247 18207
rect 22189 18167 22247 18173
rect 24489 18207 24547 18213
rect 24489 18173 24501 18207
rect 24535 18204 24547 18207
rect 24673 18207 24731 18213
rect 24673 18204 24685 18207
rect 24535 18176 24685 18204
rect 24535 18173 24547 18176
rect 24489 18167 24547 18173
rect 24673 18173 24685 18176
rect 24719 18173 24731 18207
rect 24673 18167 24731 18173
rect 24765 18207 24823 18213
rect 24765 18173 24777 18207
rect 24811 18204 24823 18207
rect 25314 18204 25320 18216
rect 24811 18176 25320 18204
rect 24811 18173 24823 18176
rect 24765 18167 24823 18173
rect 21729 18139 21787 18145
rect 21729 18105 21741 18139
rect 21775 18136 21787 18139
rect 21928 18136 21956 18167
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 25590 18164 25596 18216
rect 25648 18164 25654 18216
rect 26068 18213 26096 18244
rect 29472 18244 29929 18272
rect 25961 18207 26019 18213
rect 25961 18173 25973 18207
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 26053 18207 26111 18213
rect 26053 18173 26065 18207
rect 26099 18173 26111 18207
rect 26053 18167 26111 18173
rect 28445 18207 28503 18213
rect 28445 18173 28457 18207
rect 28491 18204 28503 18207
rect 28534 18204 28540 18216
rect 28491 18176 28540 18204
rect 28491 18173 28503 18176
rect 28445 18167 28503 18173
rect 21775 18108 21956 18136
rect 25976 18136 26004 18167
rect 28534 18164 28540 18176
rect 28592 18164 28598 18216
rect 29472 18213 29500 18244
rect 29917 18241 29929 18244
rect 29963 18241 29975 18275
rect 29917 18235 29975 18241
rect 28813 18207 28871 18213
rect 28813 18173 28825 18207
rect 28859 18204 28871 18207
rect 29089 18207 29147 18213
rect 29089 18204 29101 18207
rect 28859 18176 29101 18204
rect 28859 18173 28871 18176
rect 28813 18167 28871 18173
rect 29089 18173 29101 18176
rect 29135 18173 29147 18207
rect 29089 18167 29147 18173
rect 29181 18207 29239 18213
rect 29181 18173 29193 18207
rect 29227 18204 29239 18207
rect 29365 18207 29423 18213
rect 29365 18204 29377 18207
rect 29227 18176 29377 18204
rect 29227 18173 29239 18176
rect 29181 18167 29239 18173
rect 29365 18173 29377 18176
rect 29411 18173 29423 18207
rect 29365 18167 29423 18173
rect 29457 18207 29515 18213
rect 29457 18173 29469 18207
rect 29503 18173 29515 18207
rect 29457 18167 29515 18173
rect 29730 18164 29736 18216
rect 29788 18164 29794 18216
rect 29825 18207 29883 18213
rect 29825 18173 29837 18207
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 26145 18139 26203 18145
rect 26145 18136 26157 18139
rect 25976 18108 26157 18136
rect 21775 18105 21787 18108
rect 21729 18099 21787 18105
rect 26145 18105 26157 18108
rect 26191 18105 26203 18139
rect 26145 18099 26203 18105
rect 29641 18139 29699 18145
rect 29641 18105 29653 18139
rect 29687 18136 29699 18139
rect 29840 18136 29868 18167
rect 29687 18108 29868 18136
rect 29687 18105 29699 18108
rect 29641 18099 29699 18105
rect 22281 18071 22339 18077
rect 22281 18068 22293 18071
rect 21284 18040 22293 18068
rect 20165 18031 20223 18037
rect 22281 18037 22293 18040
rect 22327 18037 22339 18071
rect 22281 18031 22339 18037
rect 24397 18071 24455 18077
rect 24397 18037 24409 18071
rect 24443 18068 24455 18071
rect 24946 18068 24952 18080
rect 24443 18040 24952 18068
rect 24443 18037 24455 18040
rect 24397 18031 24455 18037
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25774 18028 25780 18080
rect 25832 18068 25838 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25832 18040 25881 18068
rect 25832 18028 25838 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25869 18031 25927 18037
rect 552 17978 31648 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31648 17978
rect 552 17904 31648 17926
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 2593 17867 2651 17873
rect 2593 17864 2605 17867
rect 2004 17836 2605 17864
rect 2004 17824 2010 17836
rect 2593 17833 2605 17836
rect 2639 17833 2651 17867
rect 2593 17827 2651 17833
rect 3878 17824 3884 17876
rect 3936 17824 3942 17876
rect 9674 17824 9680 17876
rect 9732 17824 9738 17876
rect 18046 17824 18052 17876
rect 18104 17824 18110 17876
rect 19061 17867 19119 17873
rect 19061 17833 19073 17867
rect 19107 17864 19119 17867
rect 19518 17864 19524 17876
rect 19107 17836 19524 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 22152 17836 22293 17864
rect 22152 17824 22158 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 25314 17824 25320 17876
rect 25372 17824 25378 17876
rect 29730 17824 29736 17876
rect 29788 17864 29794 17876
rect 30009 17867 30067 17873
rect 30009 17864 30021 17867
rect 29788 17836 30021 17864
rect 29788 17824 29794 17836
rect 30009 17833 30021 17836
rect 30055 17833 30067 17867
rect 30009 17827 30067 17833
rect 4709 17799 4767 17805
rect 4709 17796 4721 17799
rect 3988 17768 4721 17796
rect 1854 17688 1860 17740
rect 1912 17688 1918 17740
rect 1946 17688 1952 17740
rect 2004 17688 2010 17740
rect 3988 17737 4016 17768
rect 4709 17765 4721 17768
rect 4755 17765 4767 17799
rect 4709 17759 4767 17765
rect 5537 17799 5595 17805
rect 5537 17765 5549 17799
rect 5583 17796 5595 17799
rect 7101 17799 7159 17805
rect 5583 17768 5856 17796
rect 5583 17765 5595 17768
rect 5537 17759 5595 17765
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17728 2099 17731
rect 2225 17731 2283 17737
rect 2225 17728 2237 17731
rect 2087 17700 2237 17728
rect 2087 17697 2099 17700
rect 2041 17691 2099 17697
rect 2225 17697 2237 17700
rect 2271 17697 2283 17731
rect 2225 17691 2283 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2501 17731 2559 17737
rect 2501 17728 2513 17731
rect 2363 17700 2513 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2501 17697 2513 17700
rect 2547 17697 2559 17731
rect 2501 17691 2559 17697
rect 3973 17731 4031 17737
rect 3973 17697 3985 17731
rect 4019 17697 4031 17731
rect 3973 17691 4031 17697
rect 4062 17688 4068 17740
rect 4120 17688 4126 17740
rect 4157 17731 4215 17737
rect 4157 17697 4169 17731
rect 4203 17728 4215 17731
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 4203 17700 4353 17728
rect 4203 17697 4215 17700
rect 4157 17691 4215 17697
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 4341 17691 4399 17697
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 4479 17700 4629 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4617 17697 4629 17700
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 5626 17688 5632 17740
rect 5684 17688 5690 17740
rect 5828 17737 5856 17768
rect 7101 17765 7113 17799
rect 7147 17796 7159 17799
rect 12805 17799 12863 17805
rect 7147 17768 7604 17796
rect 7147 17765 7159 17768
rect 7101 17759 7159 17765
rect 5813 17731 5871 17737
rect 5813 17697 5825 17731
rect 5859 17697 5871 17731
rect 5813 17691 5871 17697
rect 5905 17731 5963 17737
rect 5905 17697 5917 17731
rect 5951 17728 5963 17731
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 5951 17700 6101 17728
rect 5951 17697 5963 17700
rect 5905 17691 5963 17697
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 6181 17731 6239 17737
rect 6181 17697 6193 17731
rect 6227 17728 6239 17731
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6227 17700 6377 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 6365 17697 6377 17700
rect 6411 17697 6423 17731
rect 6365 17691 6423 17697
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6503 17700 6745 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6871 17700 7021 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7466 17688 7472 17740
rect 7524 17688 7530 17740
rect 7576 17737 7604 17768
rect 12805 17765 12817 17799
rect 12851 17796 12863 17799
rect 13633 17799 13691 17805
rect 13633 17796 13645 17799
rect 12851 17768 13032 17796
rect 12851 17765 12863 17768
rect 12805 17759 12863 17765
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 7653 17731 7711 17737
rect 7653 17697 7665 17731
rect 7699 17728 7711 17731
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7699 17700 7941 17728
rect 7699 17697 7711 17700
rect 7653 17691 7711 17697
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 8067 17700 8217 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17728 8355 17731
rect 8481 17731 8539 17737
rect 8481 17728 8493 17731
rect 8343 17700 8493 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 8481 17697 8493 17700
rect 8527 17697 8539 17731
rect 8481 17691 8539 17697
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8757 17731 8815 17737
rect 8757 17728 8769 17731
rect 8619 17700 8769 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8757 17697 8769 17700
rect 8803 17697 8815 17731
rect 8757 17691 8815 17697
rect 8849 17731 8907 17737
rect 8849 17697 8861 17731
rect 8895 17728 8907 17731
rect 9033 17731 9091 17737
rect 9033 17728 9045 17731
rect 8895 17700 9045 17728
rect 8895 17697 8907 17700
rect 8849 17691 8907 17697
rect 9033 17697 9045 17700
rect 9079 17697 9091 17731
rect 9033 17691 9091 17697
rect 9306 17688 9312 17740
rect 9364 17688 9370 17740
rect 13004 17737 13032 17768
rect 13464 17768 13645 17796
rect 13464 17737 13492 17768
rect 13633 17765 13645 17768
rect 13679 17765 13691 17799
rect 13633 17759 13691 17765
rect 14829 17799 14887 17805
rect 14829 17765 14841 17799
rect 14875 17796 14887 17799
rect 20625 17799 20683 17805
rect 20625 17796 20637 17799
rect 14875 17768 15608 17796
rect 14875 17765 14887 17768
rect 14829 17759 14887 17765
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17697 9643 17731
rect 9585 17691 9643 17697
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17697 12679 17731
rect 12621 17691 12679 17697
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17697 12955 17731
rect 12897 17691 12955 17697
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17697 13047 17731
rect 12989 17691 13047 17697
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9600 17660 9628 17691
rect 9171 17632 9628 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 12636 17592 12664 17691
rect 12912 17660 12940 17691
rect 13538 17688 13544 17740
rect 13596 17688 13602 17740
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15580 17737 15608 17768
rect 20456 17768 20637 17796
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 15243 17700 15393 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12912 17632 13369 17660
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 15488 17660 15516 17691
rect 17586 17688 17592 17740
rect 17644 17688 17650 17740
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17819 17700 17969 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15488 17632 15669 17660
rect 13357 17623 13415 17629
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17696 17660 17724 17691
rect 18966 17688 18972 17740
rect 19024 17688 19030 17740
rect 19610 17688 19616 17740
rect 19668 17688 19674 17740
rect 20456 17737 20484 17768
rect 20625 17765 20637 17768
rect 20671 17765 20683 17799
rect 22557 17799 22615 17805
rect 22557 17796 22569 17799
rect 20625 17759 20683 17765
rect 22112 17768 22569 17796
rect 22112 17737 22140 17768
rect 22557 17765 22569 17768
rect 22603 17765 22615 17799
rect 25041 17799 25099 17805
rect 25041 17796 25053 17799
rect 22557 17759 22615 17765
rect 24872 17768 25053 17796
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19843 17700 19993 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20441 17731 20499 17737
rect 20441 17697 20453 17731
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17697 20591 17731
rect 20533 17691 20591 17697
rect 22097 17731 22155 17737
rect 22097 17697 22109 17731
rect 22143 17697 22155 17731
rect 22097 17691 22155 17697
rect 22189 17731 22247 17737
rect 22189 17697 22201 17731
rect 22235 17697 22247 17731
rect 22189 17691 22247 17697
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17728 22707 17731
rect 22833 17731 22891 17737
rect 22833 17728 22845 17731
rect 22695 17700 22845 17728
rect 22695 17697 22707 17700
rect 22649 17691 22707 17697
rect 22833 17697 22845 17700
rect 22879 17697 22891 17731
rect 22833 17691 22891 17697
rect 22925 17731 22983 17737
rect 22925 17697 22937 17731
rect 22971 17728 22983 17731
rect 23109 17731 23167 17737
rect 23109 17728 23121 17731
rect 22971 17700 23121 17728
rect 22971 17697 22983 17700
rect 22925 17691 22983 17697
rect 23109 17697 23121 17700
rect 23155 17697 23167 17731
rect 23109 17691 23167 17697
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23385 17731 23443 17737
rect 23385 17728 23397 17731
rect 23247 17700 23397 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23385 17697 23397 17700
rect 23431 17697 23443 17731
rect 23385 17691 23443 17697
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17697 23535 17731
rect 23477 17691 23535 17697
rect 17543 17632 17724 17660
rect 19521 17663 19579 17669
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 19720 17660 19748 17691
rect 19567 17632 19748 17660
rect 20073 17663 20131 17669
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20548 17660 20576 17691
rect 20119 17632 20576 17660
rect 22005 17663 22063 17669
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22204 17660 22232 17691
rect 22051 17632 22232 17660
rect 23492 17660 23520 17691
rect 23566 17688 23572 17740
rect 23624 17688 23630 17740
rect 24872 17737 24900 17768
rect 25041 17765 25053 17768
rect 25087 17765 25099 17799
rect 26789 17799 26847 17805
rect 26789 17796 26801 17799
rect 25041 17759 25099 17765
rect 26252 17768 26801 17796
rect 24029 17731 24087 17737
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24213 17731 24271 17737
rect 24213 17728 24225 17731
rect 24075 17700 24225 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 24213 17697 24225 17700
rect 24259 17697 24271 17731
rect 24213 17691 24271 17697
rect 24305 17731 24363 17737
rect 24305 17697 24317 17731
rect 24351 17728 24363 17731
rect 24489 17731 24547 17737
rect 24489 17728 24501 17731
rect 24351 17700 24501 17728
rect 24351 17697 24363 17700
rect 24305 17691 24363 17697
rect 24489 17697 24501 17700
rect 24535 17697 24547 17731
rect 24489 17691 24547 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24765 17731 24823 17737
rect 24765 17728 24777 17731
rect 24627 17700 24777 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24765 17697 24777 17700
rect 24811 17697 24823 17731
rect 24765 17691 24823 17697
rect 24857 17731 24915 17737
rect 24857 17697 24869 17731
rect 24903 17697 24915 17731
rect 24857 17691 24915 17697
rect 24946 17688 24952 17740
rect 25004 17688 25010 17740
rect 25222 17688 25228 17740
rect 25280 17688 25286 17740
rect 25774 17688 25780 17740
rect 25832 17688 25838 17740
rect 26252 17737 26280 17768
rect 26789 17765 26801 17768
rect 26835 17765 26847 17799
rect 26789 17759 26847 17765
rect 26237 17731 26295 17737
rect 26237 17697 26249 17731
rect 26283 17697 26295 17731
rect 26237 17691 26295 17697
rect 26421 17731 26479 17737
rect 26421 17697 26433 17731
rect 26467 17697 26479 17731
rect 26421 17691 26479 17697
rect 26513 17731 26571 17737
rect 26513 17697 26525 17731
rect 26559 17728 26571 17731
rect 26697 17731 26755 17737
rect 26697 17728 26709 17731
rect 26559 17700 26709 17728
rect 26559 17697 26571 17700
rect 26513 17691 26571 17697
rect 26697 17697 26709 17700
rect 26743 17697 26755 17731
rect 26697 17691 26755 17697
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23492 17632 23673 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17660 25927 17663
rect 26436 17660 26464 17691
rect 27982 17688 27988 17740
rect 28040 17728 28046 17740
rect 28077 17731 28135 17737
rect 28077 17728 28089 17731
rect 28040 17700 28089 17728
rect 28040 17688 28046 17700
rect 28077 17697 28089 17700
rect 28123 17697 28135 17731
rect 28077 17691 28135 17697
rect 29546 17688 29552 17740
rect 29604 17688 29610 17740
rect 29641 17731 29699 17737
rect 29641 17697 29653 17731
rect 29687 17697 29699 17731
rect 29641 17691 29699 17697
rect 29733 17731 29791 17737
rect 29733 17697 29745 17731
rect 29779 17728 29791 17731
rect 29917 17731 29975 17737
rect 29917 17728 29929 17731
rect 29779 17700 29929 17728
rect 29779 17697 29791 17700
rect 29733 17691 29791 17697
rect 29917 17697 29929 17700
rect 29963 17697 29975 17731
rect 29917 17691 29975 17697
rect 25915 17632 26464 17660
rect 29457 17663 29515 17669
rect 25915 17629 25927 17632
rect 25869 17623 25927 17629
rect 29457 17629 29469 17663
rect 29503 17660 29515 17663
rect 29656 17660 29684 17691
rect 29503 17632 29684 17660
rect 29503 17629 29515 17632
rect 29457 17623 29515 17629
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 12636 17564 13093 17592
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 1302 17484 1308 17536
rect 1360 17524 1366 17536
rect 1765 17527 1823 17533
rect 1765 17524 1777 17527
rect 1360 17496 1777 17524
rect 1360 17484 1366 17496
rect 1765 17493 1777 17496
rect 1811 17493 1823 17527
rect 1765 17487 1823 17493
rect 7377 17527 7435 17533
rect 7377 17493 7389 17527
rect 7423 17524 7435 17527
rect 7742 17524 7748 17536
rect 7423 17496 7748 17524
rect 7423 17493 7435 17496
rect 7377 17487 7435 17493
rect 7742 17484 7748 17496
rect 7800 17484 7806 17536
rect 9401 17527 9459 17533
rect 9401 17493 9413 17527
rect 9447 17524 9459 17527
rect 10042 17524 10048 17536
rect 9447 17496 10048 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 12529 17527 12587 17533
rect 12529 17524 12541 17527
rect 12492 17496 12541 17524
rect 12492 17484 12498 17496
rect 12529 17493 12541 17496
rect 12575 17493 12587 17527
rect 12529 17487 12587 17493
rect 15010 17484 15016 17536
rect 15068 17524 15074 17536
rect 15105 17527 15163 17533
rect 15105 17524 15117 17527
rect 15068 17496 15117 17524
rect 15068 17484 15074 17496
rect 15105 17493 15117 17496
rect 15151 17493 15163 17527
rect 15105 17487 15163 17493
rect 20254 17484 20260 17536
rect 20312 17524 20318 17536
rect 20349 17527 20407 17533
rect 20349 17524 20361 17527
rect 20312 17496 20361 17524
rect 20312 17484 20318 17496
rect 20349 17493 20361 17496
rect 20395 17493 20407 17527
rect 20349 17487 20407 17493
rect 23014 17484 23020 17536
rect 23072 17524 23078 17536
rect 23937 17527 23995 17533
rect 23937 17524 23949 17527
rect 23072 17496 23949 17524
rect 23072 17484 23078 17496
rect 23937 17493 23949 17496
rect 23983 17493 23995 17527
rect 23937 17487 23995 17493
rect 26145 17527 26203 17533
rect 26145 17493 26157 17527
rect 26191 17524 26203 17527
rect 26326 17524 26332 17536
rect 26191 17496 26332 17524
rect 26191 17493 26203 17496
rect 26145 17487 26203 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 28169 17527 28227 17533
rect 28169 17493 28181 17527
rect 28215 17524 28227 17527
rect 28994 17524 29000 17536
rect 28215 17496 29000 17524
rect 28215 17493 28227 17496
rect 28169 17487 28227 17493
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 552 17434 31648 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31648 17434
rect 552 17360 31648 17382
rect 1213 17323 1271 17329
rect 1213 17289 1225 17323
rect 1259 17320 1271 17323
rect 1946 17320 1952 17332
rect 1259 17292 1952 17320
rect 1259 17289 1271 17292
rect 1213 17283 1271 17289
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4062 17320 4068 17332
rect 4019 17292 4068 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 9033 17323 9091 17329
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9306 17320 9312 17332
rect 9079 17292 9312 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 17586 17280 17592 17332
rect 17644 17280 17650 17332
rect 22925 17323 22983 17329
rect 22925 17289 22937 17323
rect 22971 17320 22983 17323
rect 23566 17320 23572 17332
rect 22971 17292 23572 17320
rect 22971 17289 22983 17292
rect 22925 17283 22983 17289
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 25222 17320 25228 17332
rect 24903 17292 25228 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 25222 17280 25228 17292
rect 25280 17280 25286 17332
rect 29546 17280 29552 17332
rect 29604 17320 29610 17332
rect 30193 17323 30251 17329
rect 30193 17320 30205 17323
rect 29604 17292 30205 17320
rect 29604 17280 29610 17292
rect 30193 17289 30205 17292
rect 30239 17289 30251 17323
rect 30193 17283 30251 17289
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4356 17156 4813 17184
rect 1302 17076 1308 17128
rect 1360 17076 1366 17128
rect 4356 17125 4384 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 4801 17147 4859 17153
rect 7668 17156 7849 17184
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 1627 17088 1777 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1903 17088 2053 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17116 2191 17119
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 2179 17088 2329 17116
rect 2179 17085 2191 17088
rect 2133 17079 2191 17085
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17116 2467 17119
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 2455 17088 2605 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 2593 17085 2605 17088
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 2869 17119 2927 17125
rect 2869 17116 2881 17119
rect 2731 17088 2881 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 2869 17085 2881 17088
rect 2915 17085 2927 17119
rect 2869 17079 2927 17085
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3329 17119 3387 17125
rect 3329 17116 3341 17119
rect 3007 17088 3341 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3329 17085 3341 17088
rect 3375 17085 3387 17119
rect 3329 17079 3387 17085
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 3467 17088 3709 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4111 17088 4261 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 3804 17048 3832 17079
rect 4525 17051 4583 17057
rect 4525 17048 4537 17051
rect 3804 17020 4537 17048
rect 4525 17017 4537 17020
rect 4571 17017 4583 17051
rect 4632 17048 4660 17079
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 5169 17119 5227 17125
rect 5169 17085 5181 17119
rect 5215 17116 5227 17119
rect 5258 17116 5264 17128
rect 5215 17088 5264 17116
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 7668 17125 7696 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 7837 17147 7895 17153
rect 12176 17156 12633 17184
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 7742 17076 7748 17128
rect 7800 17076 7806 17128
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 9171 17088 9321 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9723 17088 9873 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 9999 17088 10149 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 10229 17119 10287 17125
rect 10229 17085 10241 17119
rect 10275 17116 10287 17119
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 10275 17088 10425 17116
rect 10275 17085 10287 17088
rect 10229 17079 10287 17085
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17116 10563 17119
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10551 17088 10701 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 10778 17076 10784 17128
rect 10836 17076 10842 17128
rect 12176 17125 12204 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 20349 17187 20407 17193
rect 14875 17156 15332 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11103 17088 11253 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 11241 17079 11299 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17116 11391 17119
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11379 17088 11529 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11609 17119 11667 17125
rect 11609 17085 11621 17119
rect 11655 17116 11667 17119
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 11655 17088 11805 17116
rect 11655 17085 11667 17088
rect 11609 17079 11667 17085
rect 11793 17085 11805 17088
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17116 11943 17119
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11931 17088 12081 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12069 17085 12081 17088
rect 12115 17085 12127 17119
rect 12069 17079 12127 17085
rect 12161 17119 12219 17125
rect 12161 17085 12173 17119
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12434 17076 12440 17128
rect 12492 17076 12498 17128
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 5077 17051 5135 17057
rect 5077 17048 5089 17051
rect 4632 17020 5089 17048
rect 4525 17011 4583 17017
rect 5077 17017 5089 17020
rect 5123 17017 5135 17051
rect 5077 17011 5135 17017
rect 12345 17051 12403 17057
rect 12345 17017 12357 17051
rect 12391 17048 12403 17051
rect 12544 17048 12572 17079
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 13688 17088 13829 17116
rect 13688 17076 13694 17088
rect 13817 17085 13829 17088
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13955 17088 14105 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14231 17088 14473 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17116 14611 17119
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14599 17088 14749 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 15010 17076 15016 17128
rect 15068 17076 15074 17128
rect 15304 17125 15332 17156
rect 20349 17153 20361 17187
rect 20395 17184 20407 17187
rect 20395 17156 20852 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 15427 17088 15761 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 15749 17085 15761 17088
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15887 17088 16037 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 16163 17088 16313 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 16301 17085 16313 17088
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17116 16451 17119
rect 16577 17119 16635 17125
rect 16577 17116 16589 17119
rect 16439 17088 16589 17116
rect 16439 17085 16451 17088
rect 16393 17079 16451 17085
rect 16577 17085 16589 17088
rect 16623 17085 16635 17119
rect 16577 17079 16635 17085
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17116 17739 17119
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17727 17088 17877 17116
rect 17727 17085 17739 17088
rect 17681 17079 17739 17085
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 18003 17088 18153 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 18279 17088 18429 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 18417 17085 18429 17088
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17116 18567 17119
rect 18785 17119 18843 17125
rect 18785 17116 18797 17119
rect 18555 17088 18797 17116
rect 18555 17085 18567 17088
rect 18509 17079 18567 17085
rect 18785 17085 18797 17088
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17116 18935 17119
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 18923 17088 19073 17116
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 12391 17020 12572 17048
rect 19168 17048 19196 17079
rect 19242 17076 19248 17128
rect 19300 17076 19306 17128
rect 20254 17076 20260 17128
rect 20312 17076 20318 17128
rect 20824 17125 20852 17156
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17085 20775 17119
rect 20717 17079 20775 17085
rect 20809 17119 20867 17125
rect 20809 17085 20821 17119
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 20901 17119 20959 17125
rect 20901 17085 20913 17119
rect 20947 17116 20959 17119
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20947 17088 21097 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 21085 17079 21143 17085
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 19168 17020 19349 17048
rect 12391 17017 12403 17020
rect 12345 17011 12403 17017
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 20732 17048 20760 17079
rect 23014 17076 23020 17128
rect 23072 17076 23078 17128
rect 24210 17076 24216 17128
rect 24268 17076 24274 17128
rect 24305 17119 24363 17125
rect 24305 17085 24317 17119
rect 24351 17116 24363 17119
rect 24489 17119 24547 17125
rect 24489 17116 24501 17119
rect 24351 17088 24501 17116
rect 24351 17085 24363 17088
rect 24305 17079 24363 17085
rect 24489 17085 24501 17088
rect 24535 17085 24547 17119
rect 24489 17079 24547 17085
rect 24581 17119 24639 17125
rect 24581 17085 24593 17119
rect 24627 17116 24639 17119
rect 24765 17119 24823 17125
rect 24765 17116 24777 17119
rect 24627 17088 24777 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 24765 17085 24777 17088
rect 24811 17085 24823 17119
rect 24765 17079 24823 17085
rect 26326 17076 26332 17128
rect 26384 17076 26390 17128
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 26605 17119 26663 17125
rect 26605 17116 26617 17119
rect 26467 17088 26617 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 26605 17085 26617 17088
rect 26651 17085 26663 17119
rect 26605 17079 26663 17085
rect 26697 17119 26755 17125
rect 26697 17085 26709 17119
rect 26743 17116 26755 17119
rect 26881 17119 26939 17125
rect 26881 17116 26893 17119
rect 26743 17088 26893 17116
rect 26743 17085 26755 17088
rect 26697 17079 26755 17085
rect 26881 17085 26893 17088
rect 26927 17085 26939 17119
rect 26881 17079 26939 17085
rect 26973 17119 27031 17125
rect 26973 17085 26985 17119
rect 27019 17116 27031 17119
rect 27157 17119 27215 17125
rect 27157 17116 27169 17119
rect 27019 17088 27169 17116
rect 27019 17085 27031 17088
rect 26973 17079 27031 17085
rect 27157 17085 27169 17088
rect 27203 17085 27215 17119
rect 27157 17079 27215 17085
rect 27249 17119 27307 17125
rect 27249 17085 27261 17119
rect 27295 17116 27307 17119
rect 27433 17119 27491 17125
rect 27433 17116 27445 17119
rect 27295 17088 27445 17116
rect 27295 17085 27307 17088
rect 27249 17079 27307 17085
rect 27433 17085 27445 17088
rect 27479 17085 27491 17119
rect 27433 17079 27491 17085
rect 27525 17119 27583 17125
rect 27525 17085 27537 17119
rect 27571 17116 27583 17119
rect 27709 17119 27767 17125
rect 27709 17116 27721 17119
rect 27571 17088 27721 17116
rect 27571 17085 27583 17088
rect 27525 17079 27583 17085
rect 27709 17085 27721 17088
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17116 27859 17119
rect 27985 17119 28043 17125
rect 27985 17116 27997 17119
rect 27847 17088 27997 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 27985 17085 27997 17088
rect 28031 17085 28043 17119
rect 27985 17079 28043 17085
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 28261 17119 28319 17125
rect 28261 17116 28273 17119
rect 28123 17088 28273 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 28261 17085 28273 17088
rect 28307 17085 28319 17119
rect 28261 17079 28319 17085
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17116 28411 17119
rect 28537 17119 28595 17125
rect 28537 17116 28549 17119
rect 28399 17088 28549 17116
rect 28399 17085 28411 17088
rect 28353 17079 28411 17085
rect 28537 17085 28549 17088
rect 28583 17085 28595 17119
rect 28537 17079 28595 17085
rect 28994 17076 29000 17128
rect 29052 17076 29058 17128
rect 29089 17119 29147 17125
rect 29089 17085 29101 17119
rect 29135 17116 29147 17119
rect 29273 17119 29331 17125
rect 29273 17116 29285 17119
rect 29135 17088 29285 17116
rect 29135 17085 29147 17088
rect 29089 17079 29147 17085
rect 29273 17085 29285 17088
rect 29319 17085 29331 17119
rect 29273 17079 29331 17085
rect 29365 17119 29423 17125
rect 29365 17085 29377 17119
rect 29411 17116 29423 17119
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 29411 17088 29561 17116
rect 29411 17085 29423 17088
rect 29365 17079 29423 17085
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 29641 17119 29699 17125
rect 29641 17085 29653 17119
rect 29687 17116 29699 17119
rect 29825 17119 29883 17125
rect 29825 17116 29837 17119
rect 29687 17088 29837 17116
rect 29687 17085 29699 17088
rect 29641 17079 29699 17085
rect 29825 17085 29837 17088
rect 29871 17085 29883 17119
rect 29825 17079 29883 17085
rect 30098 17076 30104 17128
rect 30156 17076 30162 17128
rect 21177 17051 21235 17057
rect 21177 17048 21189 17051
rect 20732 17020 21189 17048
rect 19337 17011 19395 17017
rect 21177 17017 21189 17020
rect 21223 17017 21235 17051
rect 21177 17011 21235 17017
rect 1489 16983 1547 16989
rect 1489 16949 1501 16983
rect 1535 16980 1547 16983
rect 1762 16980 1768 16992
rect 1535 16952 1768 16980
rect 1535 16949 1547 16952
rect 1489 16943 1547 16949
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 7561 16983 7619 16989
rect 7561 16949 7573 16983
rect 7607 16980 7619 16983
rect 8110 16980 8116 16992
rect 7607 16952 8116 16980
rect 7607 16949 7619 16952
rect 7561 16943 7619 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 9585 16983 9643 16989
rect 9585 16949 9597 16983
rect 9631 16980 9643 16983
rect 9766 16980 9772 16992
rect 9631 16952 9772 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10965 16983 11023 16989
rect 10965 16949 10977 16983
rect 11011 16980 11023 16983
rect 11146 16980 11152 16992
rect 11011 16952 11152 16980
rect 11011 16949 11023 16952
rect 10965 16943 11023 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 15105 16983 15163 16989
rect 15105 16949 15117 16983
rect 15151 16980 15163 16983
rect 15378 16980 15384 16992
rect 15151 16952 15384 16980
rect 15151 16949 15163 16952
rect 15105 16943 15163 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 20625 16983 20683 16989
rect 20625 16949 20637 16983
rect 20671 16980 20683 16983
rect 20714 16980 20720 16992
rect 20671 16952 20720 16980
rect 20671 16949 20683 16952
rect 20625 16943 20683 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 28074 16940 28080 16992
rect 28132 16980 28138 16992
rect 28629 16983 28687 16989
rect 28629 16980 28641 16983
rect 28132 16952 28641 16980
rect 28132 16940 28138 16952
rect 28629 16949 28641 16952
rect 28675 16949 28687 16983
rect 28629 16943 28687 16949
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 29917 16983 29975 16989
rect 29917 16980 29929 16983
rect 29420 16952 29929 16980
rect 29420 16940 29426 16952
rect 29917 16949 29929 16952
rect 29963 16949 29975 16983
rect 29917 16943 29975 16949
rect 552 16890 31648 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31648 16890
rect 552 16816 31648 16838
rect 1854 16736 1860 16788
rect 1912 16736 1918 16788
rect 4890 16736 4896 16788
rect 4948 16736 4954 16788
rect 5258 16736 5264 16788
rect 5316 16736 5322 16788
rect 9398 16736 9404 16788
rect 9456 16776 9462 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9456 16748 9873 16776
rect 9456 16736 9462 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 11241 16779 11299 16785
rect 11241 16776 11253 16779
rect 10836 16748 11253 16776
rect 10836 16736 10842 16748
rect 11241 16745 11253 16748
rect 11287 16745 11299 16779
rect 11241 16739 11299 16745
rect 13630 16736 13636 16788
rect 13688 16736 13694 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 19242 16776 19248 16788
rect 18831 16748 19248 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 24489 16779 24547 16785
rect 24489 16776 24501 16779
rect 24044 16748 24501 16776
rect 6457 16711 6515 16717
rect 6457 16708 6469 16711
rect 6012 16680 6469 16708
rect 1762 16600 1768 16652
rect 1820 16600 1826 16652
rect 4246 16600 4252 16652
rect 4304 16600 4310 16652
rect 6012 16649 6040 16680
rect 6457 16677 6469 16680
rect 6503 16677 6515 16711
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 6457 16671 6515 16677
rect 8036 16680 8217 16708
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 4387 16612 4537 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16640 4675 16643
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4663 16612 4813 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5537 16643 5595 16649
rect 5537 16640 5549 16643
rect 5399 16612 5549 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5537 16609 5549 16612
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 5905 16643 5963 16649
rect 5905 16640 5917 16643
rect 5675 16612 5917 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5905 16609 5917 16612
rect 5951 16609 5963 16643
rect 5905 16603 5963 16609
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 6086 16600 6092 16652
rect 6144 16600 6150 16652
rect 8036 16649 8064 16680
rect 8205 16677 8217 16680
rect 8251 16677 8263 16711
rect 10137 16711 10195 16717
rect 10137 16708 10149 16711
rect 8205 16671 8263 16677
rect 9600 16680 10149 16708
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 6227 16612 6377 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6365 16609 6377 16612
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 7929 16643 7987 16649
rect 7929 16640 7941 16643
rect 7791 16612 7941 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 7929 16609 7941 16612
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 9600 16649 9628 16680
rect 10137 16677 10149 16680
rect 10183 16677 10195 16711
rect 14185 16711 14243 16717
rect 14185 16708 14197 16711
rect 10137 16671 10195 16677
rect 14016 16680 14197 16708
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9355 16612 9505 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9766 16600 9772 16652
rect 9824 16600 9830 16652
rect 10042 16600 10048 16652
rect 10100 16600 10106 16652
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 13170 16600 13176 16652
rect 13228 16600 13234 16652
rect 14016 16649 14044 16680
rect 14185 16677 14197 16680
rect 14231 16677 14243 16711
rect 15473 16711 15531 16717
rect 15473 16708 15485 16711
rect 14185 16671 14243 16677
rect 15304 16680 15485 16708
rect 15304 16649 15332 16680
rect 15473 16677 15485 16680
rect 15519 16677 15531 16711
rect 17313 16711 17371 16717
rect 17313 16708 17325 16711
rect 15473 16671 15531 16677
rect 17144 16680 17325 16708
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13725 16643 13783 16649
rect 13311 16612 13584 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13556 16572 13584 16612
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13771 16612 13921 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16609 14059 16643
rect 14001 16603 14059 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 14108 16572 14136 16603
rect 15378 16600 15384 16652
rect 15436 16600 15442 16652
rect 16666 16600 16672 16652
rect 16724 16600 16730 16652
rect 17144 16649 17172 16680
rect 17313 16677 17325 16680
rect 17359 16677 17371 16711
rect 19613 16711 19671 16717
rect 19613 16708 19625 16711
rect 17313 16671 17371 16677
rect 18892 16680 19625 16708
rect 18892 16649 18920 16680
rect 19613 16677 19625 16680
rect 19659 16677 19671 16711
rect 19613 16671 19671 16677
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17129 16643 17187 16649
rect 16807 16612 17080 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 13556 16544 14136 16572
rect 17052 16572 17080 16612
rect 17129 16609 17141 16643
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16609 18935 16643
rect 18877 16603 18935 16609
rect 17236 16572 17264 16603
rect 18966 16600 18972 16652
rect 19024 16600 19030 16652
rect 19061 16643 19119 16649
rect 19061 16609 19073 16643
rect 19107 16640 19119 16643
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 19107 16612 19257 16640
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 19245 16609 19257 16612
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16640 19395 16643
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 19383 16612 19533 16640
rect 19383 16609 19395 16612
rect 19337 16603 19395 16609
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 20714 16600 20720 16652
rect 20772 16600 20778 16652
rect 24044 16649 24072 16748
rect 24489 16745 24501 16748
rect 24535 16745 24547 16779
rect 24489 16739 24547 16745
rect 27982 16736 27988 16788
rect 28040 16736 28046 16788
rect 29273 16779 29331 16785
rect 29273 16745 29285 16779
rect 29319 16776 29331 16779
rect 30098 16776 30104 16788
rect 29319 16748 30104 16776
rect 29319 16745 29331 16748
rect 29273 16739 29331 16745
rect 30098 16736 30104 16748
rect 30156 16736 30162 16788
rect 24213 16711 24271 16717
rect 24213 16677 24225 16711
rect 24259 16708 24271 16711
rect 25041 16711 25099 16717
rect 25041 16708 25053 16711
rect 24259 16680 24440 16708
rect 24259 16677 24271 16680
rect 24213 16671 24271 16677
rect 24412 16649 24440 16680
rect 24872 16680 25053 16708
rect 24872 16649 24900 16680
rect 25041 16677 25053 16680
rect 25087 16677 25099 16711
rect 25041 16671 25099 16677
rect 29825 16711 29883 16717
rect 29825 16677 29837 16711
rect 29871 16708 29883 16711
rect 30374 16708 30380 16720
rect 29871 16680 30380 16708
rect 29871 16677 29883 16680
rect 29825 16671 29883 16677
rect 30374 16668 30380 16680
rect 30432 16668 30438 16720
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16640 20867 16643
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20855 16612 21281 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21361 16643 21419 16649
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21407 16612 21557 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 21545 16603 21603 16609
rect 21637 16643 21695 16649
rect 21637 16609 21649 16643
rect 21683 16640 21695 16643
rect 21821 16643 21879 16649
rect 21821 16640 21833 16643
rect 21683 16612 21833 16640
rect 21683 16609 21695 16612
rect 21637 16603 21695 16609
rect 21821 16609 21833 16612
rect 21867 16609 21879 16643
rect 21821 16603 21879 16609
rect 21913 16643 21971 16649
rect 21913 16609 21925 16643
rect 21959 16640 21971 16643
rect 22097 16643 22155 16649
rect 22097 16640 22109 16643
rect 21959 16612 22109 16640
rect 21959 16609 21971 16612
rect 21913 16603 21971 16609
rect 22097 16609 22109 16612
rect 22143 16609 22155 16643
rect 22097 16603 22155 16609
rect 22189 16643 22247 16649
rect 22189 16609 22201 16643
rect 22235 16640 22247 16643
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22235 16612 22385 16640
rect 22235 16609 22247 16612
rect 22189 16603 22247 16609
rect 22373 16609 22385 16612
rect 22419 16609 22431 16643
rect 22373 16603 22431 16609
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16640 22523 16643
rect 22649 16643 22707 16649
rect 22649 16640 22661 16643
rect 22511 16612 22661 16640
rect 22511 16609 22523 16612
rect 22465 16603 22523 16609
rect 22649 16609 22661 16612
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16609 24087 16643
rect 24029 16603 24087 16609
rect 24305 16643 24363 16649
rect 24305 16609 24317 16643
rect 24351 16609 24363 16643
rect 24305 16603 24363 16609
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16609 24455 16643
rect 24765 16643 24823 16649
rect 24765 16640 24777 16643
rect 24397 16603 24455 16609
rect 24596 16612 24777 16640
rect 17052 16544 17264 16572
rect 24320 16572 24348 16603
rect 24596 16572 24624 16612
rect 24765 16609 24777 16612
rect 24811 16609 24823 16643
rect 24765 16603 24823 16609
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 24946 16600 24952 16652
rect 25004 16600 25010 16652
rect 25501 16643 25559 16649
rect 25501 16609 25513 16643
rect 25547 16640 25559 16643
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 25547 16612 25697 16640
rect 25547 16609 25559 16612
rect 25501 16603 25559 16609
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 25961 16643 26019 16649
rect 25961 16640 25973 16643
rect 25823 16612 25973 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 25961 16609 25973 16612
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26050 16600 26056 16652
rect 26108 16600 26114 16652
rect 28074 16600 28080 16652
rect 28132 16600 28138 16652
rect 29362 16600 29368 16652
rect 29420 16600 29426 16652
rect 29914 16600 29920 16652
rect 29972 16600 29978 16652
rect 24320 16544 24624 16572
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7432 16408 7665 16436
rect 7432 16396 7438 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7653 16399 7711 16405
rect 9217 16439 9275 16445
rect 9217 16405 9229 16439
rect 9263 16436 9275 16439
rect 9582 16436 9588 16448
rect 9263 16408 9588 16436
rect 9263 16405 9275 16408
rect 9217 16399 9275 16405
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 15194 16396 15200 16448
rect 15252 16396 15258 16448
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 17037 16439 17095 16445
rect 17037 16436 17049 16439
rect 17000 16408 17049 16436
rect 17000 16396 17006 16408
rect 17037 16405 17049 16408
rect 17083 16405 17095 16439
rect 17037 16399 17095 16405
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 22244 16408 22753 16436
rect 22244 16396 22250 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 23937 16439 23995 16445
rect 23937 16405 23949 16439
rect 23983 16436 23995 16439
rect 24118 16436 24124 16448
rect 23983 16408 24124 16436
rect 23983 16405 23995 16408
rect 23937 16399 23995 16405
rect 24118 16396 24124 16408
rect 24176 16396 24182 16448
rect 25406 16396 25412 16448
rect 25464 16396 25470 16448
rect 552 16346 31648 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31648 16346
rect 552 16272 31648 16294
rect 3881 16235 3939 16241
rect 3881 16201 3893 16235
rect 3927 16232 3939 16235
rect 4246 16232 4252 16244
rect 3927 16204 4252 16232
rect 3927 16201 3939 16204
rect 3881 16195 3939 16201
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6144 16204 6193 16232
rect 6144 16192 6150 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 12805 16235 12863 16241
rect 12805 16201 12817 16235
rect 12851 16232 12863 16235
rect 13170 16232 13176 16244
rect 12851 16204 13176 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 18877 16235 18935 16241
rect 18877 16201 18889 16235
rect 18923 16232 18935 16235
rect 18966 16232 18972 16244
rect 18923 16204 18972 16232
rect 18923 16201 18935 16204
rect 18877 16195 18935 16201
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 24210 16192 24216 16244
rect 24268 16192 24274 16244
rect 24765 16235 24823 16241
rect 24765 16201 24777 16235
rect 24811 16232 24823 16235
rect 24946 16232 24952 16244
rect 24811 16204 24952 16232
rect 24811 16201 24823 16204
rect 24765 16195 24823 16201
rect 24946 16192 24952 16204
rect 25004 16192 25010 16244
rect 25961 16235 26019 16241
rect 25961 16201 25973 16235
rect 26007 16232 26019 16235
rect 26050 16232 26056 16244
rect 26007 16204 26056 16232
rect 26007 16201 26019 16204
rect 25961 16195 26019 16201
rect 26050 16192 26056 16204
rect 26108 16192 26114 16244
rect 29914 16192 29920 16244
rect 29972 16232 29978 16244
rect 30193 16235 30251 16241
rect 30193 16232 30205 16235
rect 29972 16204 30205 16232
rect 29972 16192 29978 16204
rect 30193 16201 30205 16204
rect 30239 16201 30251 16235
rect 30193 16195 30251 16201
rect 4798 16096 4804 16108
rect 4540 16068 4804 16096
rect 4540 16037 4568 16068
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 6457 16099 6515 16105
rect 6457 16065 6469 16099
rect 6503 16096 6515 16099
rect 7285 16099 7343 16105
rect 6503 16068 6684 16096
rect 6503 16065 6515 16068
rect 6457 16059 6515 16065
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 16028 4307 16031
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 4295 16000 4445 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 16028 4767 16031
rect 4893 16031 4951 16037
rect 4893 16028 4905 16031
rect 4755 16000 4905 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 4893 15997 4905 16000
rect 4939 15997 4951 16031
rect 4893 15991 4951 15997
rect 6273 16031 6331 16037
rect 6273 15997 6285 16031
rect 6319 15997 6331 16031
rect 6273 15991 6331 15997
rect 3988 15892 4016 15991
rect 4157 15963 4215 15969
rect 4157 15929 4169 15963
rect 4203 15960 4215 15963
rect 4632 15960 4660 15991
rect 4203 15932 4660 15960
rect 6288 15960 6316 15991
rect 6546 15988 6552 16040
rect 6604 15988 6610 16040
rect 6656 16037 6684 16068
rect 7285 16065 7297 16099
rect 7331 16096 7343 16099
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 7331 16068 7512 16096
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 16028 6791 16031
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6779 16000 6929 16028
rect 6779 15997 6791 16000
rect 6733 15991 6791 15997
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 7374 15988 7380 16040
rect 7432 15988 7438 16040
rect 7484 16037 7512 16068
rect 9232 16068 9689 16096
rect 9232 16037 9260 16068
rect 9677 16065 9689 16068
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 11195 16068 11744 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 7561 16031 7619 16037
rect 7561 15997 7573 16031
rect 7607 16028 7619 16031
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7607 16000 7757 16028
rect 7607 15997 7619 16000
rect 7561 15991 7619 15997
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 16028 7895 16031
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7883 16000 8033 16028
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 8159 16000 8401 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 16028 8539 16031
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8527 16000 8677 16028
rect 8527 15997 8539 16000
rect 8481 15991 8539 15997
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 7009 15963 7067 15969
rect 7009 15960 7021 15963
rect 6288 15932 7021 15960
rect 4203 15929 4215 15932
rect 4157 15923 4215 15929
rect 7009 15929 7021 15932
rect 7055 15929 7067 15963
rect 7009 15923 7067 15929
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 9324 15960 9352 15991
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11716 16037 11744 16068
rect 12912 16068 13921 16096
rect 12912 16037 12940 16068
rect 13909 16065 13921 16068
rect 13955 16065 13967 16099
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 13909 16059 13967 16065
rect 15764 16068 15945 16096
rect 11609 16031 11667 16037
rect 11609 15997 11621 16031
rect 11655 15997 11667 16031
rect 11609 15991 11667 15997
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 8803 15932 9352 15960
rect 11624 15960 11652 15991
rect 13170 15988 13176 16040
rect 13228 15988 13234 16040
rect 13541 16031 13599 16037
rect 13541 15997 13553 16031
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13679 16000 13829 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 16028 14979 16031
rect 15102 16028 15108 16040
rect 14967 16000 15108 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 11793 15963 11851 15969
rect 11793 15960 11805 15963
rect 11624 15932 11805 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 11793 15929 11805 15932
rect 11839 15929 11851 15963
rect 11793 15923 11851 15929
rect 13081 15963 13139 15969
rect 13081 15929 13093 15963
rect 13127 15960 13139 15963
rect 13556 15960 13584 15991
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15764 16037 15792 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 15933 16059 15991 16065
rect 17512 16068 17693 16096
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 16028 15255 16031
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 15243 16000 15393 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 15381 15991 15439 15997
rect 15473 16031 15531 16037
rect 15473 15997 15485 16031
rect 15519 16028 15531 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15519 16000 15669 16028
rect 15519 15997 15531 16000
rect 15473 15991 15531 15997
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 15997 15899 16031
rect 15841 15991 15899 15997
rect 13127 15932 13584 15960
rect 14829 15963 14887 15969
rect 13127 15929 13139 15932
rect 13081 15923 13139 15929
rect 14829 15929 14841 15963
rect 14875 15960 14887 15963
rect 15856 15960 15884 15991
rect 16942 15988 16948 16040
rect 17000 15988 17006 16040
rect 17512 16037 17540 16068
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 19153 16099 19211 16105
rect 19153 16065 19165 16099
rect 19199 16096 19211 16099
rect 22097 16099 22155 16105
rect 19199 16068 19380 16096
rect 19199 16065 19211 16068
rect 19153 16059 19211 16065
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 17267 16000 17417 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17405 15997 17417 16000
rect 17451 15997 17463 16031
rect 17405 15991 17463 15997
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 15997 17647 16031
rect 17589 15991 17647 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 14875 15932 15884 15960
rect 16853 15963 16911 15969
rect 14875 15929 14887 15932
rect 14829 15923 14887 15929
rect 16853 15929 16865 15963
rect 16899 15960 16911 15963
rect 17604 15960 17632 15991
rect 16899 15932 17632 15960
rect 18984 15960 19012 15991
rect 19242 15988 19248 16040
rect 19300 15988 19306 16040
rect 19352 16037 19380 16068
rect 22097 16065 22109 16099
rect 22143 16096 22155 16099
rect 22143 16068 22324 16096
rect 22143 16065 22155 16068
rect 22097 16059 22155 16065
rect 19337 16031 19395 16037
rect 19337 15997 19349 16031
rect 19383 15997 19395 16031
rect 19337 15991 19395 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 19475 16000 19625 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 22186 15988 22192 16040
rect 22244 15988 22250 16040
rect 22296 16037 22324 16068
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 16028 22431 16031
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22419 16000 22569 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 16028 22707 16031
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22695 16000 22845 16028
rect 22695 15997 22707 16000
rect 22649 15991 22707 15997
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 16028 22983 16031
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 22971 16000 23121 16028
rect 22971 15997 22983 16000
rect 22925 15991 22983 15997
rect 23109 15997 23121 16000
rect 23155 15997 23167 16031
rect 23109 15991 23167 15997
rect 23201 16031 23259 16037
rect 23201 15997 23213 16031
rect 23247 16028 23259 16031
rect 23385 16031 23443 16037
rect 23385 16028 23397 16031
rect 23247 16000 23397 16028
rect 23247 15997 23259 16000
rect 23201 15991 23259 15997
rect 23385 15997 23397 16000
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 16028 24915 16031
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 24903 16000 25053 16028
rect 24903 15997 24915 16000
rect 24857 15991 24915 15997
rect 25041 15997 25053 16000
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 25133 16031 25191 16037
rect 25133 15997 25145 16031
rect 25179 16028 25191 16031
rect 25317 16031 25375 16037
rect 25317 16028 25329 16031
rect 25179 16000 25329 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 25317 15997 25329 16000
rect 25363 15997 25375 16031
rect 25317 15991 25375 15997
rect 25406 15988 25412 16040
rect 25464 15988 25470 16040
rect 26053 16031 26111 16037
rect 26053 15997 26065 16031
rect 26099 16028 26111 16031
rect 26237 16031 26295 16037
rect 26237 16028 26249 16031
rect 26099 16000 26249 16028
rect 26099 15997 26111 16000
rect 26053 15991 26111 15997
rect 26237 15997 26249 16000
rect 26283 15997 26295 16031
rect 26237 15991 26295 15997
rect 26329 16031 26387 16037
rect 26329 15997 26341 16031
rect 26375 16028 26387 16031
rect 26513 16031 26571 16037
rect 26513 16028 26525 16031
rect 26375 16000 26525 16028
rect 26375 15997 26387 16000
rect 26329 15991 26387 15997
rect 26513 15997 26525 16000
rect 26559 15997 26571 16031
rect 26513 15991 26571 15997
rect 26605 16031 26663 16037
rect 26605 15997 26617 16031
rect 26651 16028 26663 16031
rect 26789 16031 26847 16037
rect 26789 16028 26801 16031
rect 26651 16000 26801 16028
rect 26651 15997 26663 16000
rect 26605 15991 26663 15997
rect 26789 15997 26801 16000
rect 26835 15997 26847 16031
rect 26789 15991 26847 15997
rect 26881 16031 26939 16037
rect 26881 15997 26893 16031
rect 26927 16028 26939 16031
rect 27065 16031 27123 16037
rect 27065 16028 27077 16031
rect 26927 16000 27077 16028
rect 26927 15997 26939 16000
rect 26881 15991 26939 15997
rect 27065 15997 27077 16000
rect 27111 15997 27123 16031
rect 27065 15991 27123 15997
rect 27157 16031 27215 16037
rect 27157 15997 27169 16031
rect 27203 16028 27215 16031
rect 27341 16031 27399 16037
rect 27341 16028 27353 16031
rect 27203 16000 27353 16028
rect 27203 15997 27215 16000
rect 27157 15991 27215 15997
rect 27341 15997 27353 16000
rect 27387 15997 27399 16031
rect 27341 15991 27399 15997
rect 27433 16031 27491 16037
rect 27433 15997 27445 16031
rect 27479 16028 27491 16031
rect 27617 16031 27675 16037
rect 27617 16028 27629 16031
rect 27479 16000 27629 16028
rect 27479 15997 27491 16000
rect 27433 15991 27491 15997
rect 27617 15997 27629 16000
rect 27663 15997 27675 16031
rect 27617 15991 27675 15997
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 27893 16031 27951 16037
rect 27893 16028 27905 16031
rect 27755 16000 27905 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 27893 15997 27905 16000
rect 27939 15997 27951 16031
rect 27893 15991 27951 15997
rect 27985 16031 28043 16037
rect 27985 15997 27997 16031
rect 28031 16028 28043 16031
rect 28169 16031 28227 16037
rect 28169 16028 28181 16031
rect 28031 16000 28181 16028
rect 28031 15997 28043 16000
rect 27985 15991 28043 15997
rect 28169 15997 28181 16000
rect 28215 15997 28227 16031
rect 28169 15991 28227 15997
rect 28261 16031 28319 16037
rect 28261 15997 28273 16031
rect 28307 16028 28319 16031
rect 28445 16031 28503 16037
rect 28445 16028 28457 16031
rect 28307 16000 28457 16028
rect 28307 15997 28319 16000
rect 28261 15991 28319 15997
rect 28445 15997 28457 16000
rect 28491 15997 28503 16031
rect 28445 15991 28503 15997
rect 28537 16031 28595 16037
rect 28537 15997 28549 16031
rect 28583 16028 28595 16031
rect 28721 16031 28779 16037
rect 28721 16028 28733 16031
rect 28583 16000 28733 16028
rect 28583 15997 28595 16000
rect 28537 15991 28595 15997
rect 28721 15997 28733 16000
rect 28767 15997 28779 16031
rect 28721 15991 28779 15997
rect 28813 16031 28871 16037
rect 28813 15997 28825 16031
rect 28859 16028 28871 16031
rect 29089 16031 29147 16037
rect 29089 16028 29101 16031
rect 28859 16000 29101 16028
rect 28859 15997 28871 16000
rect 28813 15991 28871 15997
rect 29089 15997 29101 16000
rect 29135 15997 29147 16031
rect 29089 15991 29147 15997
rect 29181 16031 29239 16037
rect 29181 15997 29193 16031
rect 29227 16028 29239 16031
rect 29365 16031 29423 16037
rect 29365 16028 29377 16031
rect 29227 16000 29377 16028
rect 29227 15997 29239 16000
rect 29181 15991 29239 15997
rect 29365 15997 29377 16000
rect 29411 15997 29423 16031
rect 29365 15991 29423 15997
rect 29457 16031 29515 16037
rect 29457 15997 29469 16031
rect 29503 16028 29515 16031
rect 29641 16031 29699 16037
rect 29641 16028 29653 16031
rect 29503 16000 29653 16028
rect 29503 15997 29515 16000
rect 29457 15991 29515 15997
rect 29641 15997 29653 16000
rect 29687 15997 29699 16031
rect 29641 15991 29699 15997
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 29917 16031 29975 16037
rect 29917 16028 29929 16031
rect 29779 16000 29929 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 29917 15997 29929 16000
rect 29963 15997 29975 16031
rect 29917 15991 29975 15997
rect 30009 16031 30067 16037
rect 30009 15997 30021 16031
rect 30055 15997 30067 16031
rect 30009 15991 30067 15997
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 18984 15932 19717 15960
rect 16899 15929 16911 15932
rect 16853 15923 16911 15929
rect 19705 15929 19717 15932
rect 19751 15929 19763 15963
rect 30024 15960 30052 15991
rect 30098 15988 30104 16040
rect 30156 15988 30162 16040
rect 30374 15988 30380 16040
rect 30432 15988 30438 16040
rect 30469 15963 30527 15969
rect 30469 15960 30481 15963
rect 30024 15932 30481 15960
rect 19705 15923 19763 15929
rect 30469 15929 30481 15932
rect 30515 15929 30527 15963
rect 30469 15923 30527 15929
rect 4985 15895 5043 15901
rect 4985 15892 4997 15895
rect 3988 15864 4997 15892
rect 4985 15861 4997 15864
rect 5031 15861 5043 15895
rect 4985 15855 5043 15861
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8996 15864 9137 15892
rect 8996 15852 9002 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 9398 15852 9404 15904
rect 9456 15852 9462 15904
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 11606 15892 11612 15904
rect 11563 15864 11612 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15746 15892 15752 15904
rect 15151 15864 15752 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17586 15892 17592 15904
rect 17175 15864 17592 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23477 15895 23535 15901
rect 23477 15892 23489 15895
rect 23164 15864 23489 15892
rect 23164 15852 23170 15864
rect 23477 15861 23489 15864
rect 23523 15861 23535 15895
rect 23477 15855 23535 15861
rect 552 15802 31648 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31648 15802
rect 552 15728 31648 15750
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 4893 15691 4951 15697
rect 4893 15688 4905 15691
rect 4856 15660 4905 15688
rect 4856 15648 4862 15660
rect 4893 15657 4905 15660
rect 4939 15657 4951 15691
rect 4893 15651 4951 15657
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6604 15660 6929 15688
rect 6604 15648 6610 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 13170 15648 13176 15700
rect 13228 15648 13234 15700
rect 19242 15648 19248 15700
rect 19300 15688 19306 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19300 15660 19809 15688
rect 19300 15648 19306 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 19797 15651 19855 15657
rect 30098 15648 30104 15700
rect 30156 15648 30162 15700
rect 11333 15623 11391 15629
rect 11333 15620 11345 15623
rect 11164 15592 11345 15620
rect 3970 15512 3976 15564
rect 4028 15512 4034 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4249 15555 4307 15561
rect 4249 15552 4261 15555
rect 4111 15524 4261 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4249 15521 4261 15524
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 4387 15524 4537 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4663 15524 4813 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15552 6423 15555
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 6411 15524 6561 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6687 15524 6837 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 8938 15512 8944 15564
rect 8996 15512 9002 15564
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 8849 15487 8907 15493
rect 8849 15453 8861 15487
rect 8895 15484 8907 15487
rect 9048 15484 9076 15515
rect 9398 15512 9404 15564
rect 9456 15512 9462 15564
rect 11164 15561 11192 15592
rect 11333 15589 11345 15592
rect 11379 15589 11391 15623
rect 11333 15583 11391 15589
rect 12897 15623 12955 15629
rect 12897 15589 12909 15623
rect 12943 15620 12955 15623
rect 19610 15620 19616 15632
rect 12943 15592 13124 15620
rect 12943 15589 12955 15592
rect 12897 15583 12955 15589
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15552 9551 15555
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9539 15524 9781 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9907 15524 10057 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10183 15524 10333 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10459 15524 10609 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 8895 15456 9076 15484
rect 10689 15487 10747 15493
rect 8895 15453 8907 15456
rect 8849 15447 8907 15453
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 11256 15484 11284 15515
rect 11606 15512 11612 15564
rect 11664 15512 11670 15564
rect 13096 15561 13124 15592
rect 19076 15592 19616 15620
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15552 11759 15555
rect 11885 15555 11943 15561
rect 11885 15552 11897 15555
rect 11747 15524 11897 15552
rect 11747 15521 11759 15524
rect 11701 15515 11759 15521
rect 11885 15521 11897 15524
rect 11931 15521 11943 15555
rect 11885 15515 11943 15521
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 12023 15524 12173 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12437 15555 12495 15561
rect 12437 15552 12449 15555
rect 12299 15524 12449 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12437 15521 12449 15524
rect 12483 15521 12495 15555
rect 12437 15515 12495 15521
rect 12989 15555 13047 15561
rect 12989 15521 13001 15555
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14829 15555 14887 15561
rect 13403 15524 13584 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 10735 15456 11284 15484
rect 13004 15484 13032 15515
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13004 15456 13461 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 12529 15419 12587 15425
rect 12529 15385 12541 15419
rect 12575 15416 12587 15419
rect 13556 15416 13584 15524
rect 14829 15521 14841 15555
rect 14875 15552 14887 15555
rect 15013 15555 15071 15561
rect 15013 15552 15025 15555
rect 14875 15524 15025 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 15013 15521 15025 15524
rect 15059 15521 15071 15555
rect 15013 15515 15071 15521
rect 15105 15555 15163 15561
rect 15105 15521 15117 15555
rect 15151 15552 15163 15555
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15151 15524 15301 15552
rect 15151 15521 15163 15524
rect 15105 15515 15163 15521
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 15427 15524 15577 15552
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 15672 15484 15700 15515
rect 15746 15512 15752 15564
rect 15804 15512 15810 15564
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15552 17003 15555
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 16991 15524 17141 15552
rect 16991 15521 17003 15524
rect 16945 15515 17003 15521
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 17405 15555 17463 15561
rect 17405 15552 17417 15555
rect 17267 15524 17417 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 17405 15521 17417 15524
rect 17451 15521 17463 15555
rect 17405 15515 17463 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15672 15456 15853 15484
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 17512 15484 17540 15515
rect 17586 15512 17592 15564
rect 17644 15512 17650 15564
rect 19076 15561 19104 15592
rect 19610 15580 19616 15592
rect 19668 15580 19674 15632
rect 23569 15623 23627 15629
rect 23569 15589 23581 15623
rect 23615 15620 23627 15623
rect 29273 15623 29331 15629
rect 23615 15592 24072 15620
rect 23615 15589 23627 15592
rect 23569 15583 23627 15589
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 19153 15555 19211 15561
rect 19153 15521 19165 15555
rect 19199 15521 19211 15555
rect 19153 15515 19211 15521
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15552 19303 15555
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19291 15524 19441 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 19567 15524 19717 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 19705 15521 19717 15524
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17512 15456 17693 15484
rect 15841 15447 15899 15453
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19168 15484 19196 15515
rect 22094 15512 22100 15564
rect 22152 15512 22158 15564
rect 23106 15512 23112 15564
rect 23164 15512 23170 15564
rect 24044 15561 24072 15592
rect 29273 15589 29285 15623
rect 29319 15620 29331 15623
rect 29319 15592 29500 15620
rect 29319 15589 29331 15592
rect 29273 15583 29331 15589
rect 23201 15555 23259 15561
rect 23201 15521 23213 15555
rect 23247 15521 23259 15555
rect 23201 15515 23259 15521
rect 23293 15555 23351 15561
rect 23293 15521 23305 15555
rect 23339 15552 23351 15555
rect 23477 15555 23535 15561
rect 23477 15552 23489 15555
rect 23339 15524 23489 15552
rect 23339 15521 23351 15524
rect 23293 15515 23351 15521
rect 23477 15521 23489 15524
rect 23523 15521 23535 15555
rect 23477 15515 23535 15521
rect 23937 15555 23995 15561
rect 23937 15521 23949 15555
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 24029 15555 24087 15561
rect 24029 15521 24041 15555
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 24305 15555 24363 15561
rect 24305 15521 24317 15555
rect 24351 15521 24363 15555
rect 24305 15515 24363 15521
rect 19015 15456 19196 15484
rect 23017 15487 23075 15493
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 23017 15453 23029 15487
rect 23063 15484 23075 15487
rect 23216 15484 23244 15515
rect 23063 15456 23244 15484
rect 23952 15484 23980 15515
rect 24121 15487 24179 15493
rect 24121 15484 24133 15487
rect 23952 15456 24133 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 24121 15453 24133 15456
rect 24167 15453 24179 15487
rect 24121 15447 24179 15453
rect 12575 15388 13584 15416
rect 23845 15419 23903 15425
rect 12575 15385 12587 15388
rect 12529 15379 12587 15385
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24320 15416 24348 15515
rect 29362 15512 29368 15564
rect 29420 15512 29426 15564
rect 29472 15561 29500 15592
rect 29457 15555 29515 15561
rect 29457 15521 29469 15555
rect 29503 15521 29515 15555
rect 29457 15515 29515 15521
rect 29549 15555 29607 15561
rect 29549 15521 29561 15555
rect 29595 15552 29607 15555
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 29595 15524 29745 15552
rect 29595 15521 29607 15524
rect 29549 15515 29607 15521
rect 29733 15521 29745 15524
rect 29779 15521 29791 15555
rect 29733 15515 29791 15521
rect 29825 15555 29883 15561
rect 29825 15521 29837 15555
rect 29871 15552 29883 15555
rect 30009 15555 30067 15561
rect 30009 15552 30021 15555
rect 29871 15524 30021 15552
rect 29871 15521 29883 15524
rect 29825 15515 29883 15521
rect 30009 15521 30021 15524
rect 30055 15521 30067 15555
rect 30009 15515 30067 15521
rect 23891 15388 24348 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 14826 15348 14832 15360
rect 14783 15320 14832 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 16853 15351 16911 15357
rect 16853 15317 16865 15351
rect 16899 15348 16911 15351
rect 17218 15348 17224 15360
rect 16899 15320 17224 15348
rect 16899 15317 16911 15320
rect 16853 15311 16911 15317
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15348 22247 15351
rect 22738 15348 22744 15360
rect 22235 15320 22744 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 22738 15308 22744 15320
rect 22796 15308 22802 15360
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 24397 15351 24455 15357
rect 24397 15348 24409 15351
rect 23716 15320 24409 15348
rect 23716 15308 23722 15320
rect 24397 15317 24409 15320
rect 24443 15317 24455 15351
rect 24397 15311 24455 15317
rect 552 15258 31648 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31648 15258
rect 552 15184 31648 15206
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4062 15144 4068 15156
rect 3835 15116 4068 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 6270 15144 6276 15156
rect 6043 15116 6276 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 19610 15104 19616 15156
rect 19668 15104 19674 15156
rect 29362 15104 29368 15156
rect 29420 15144 29426 15156
rect 29917 15147 29975 15153
rect 29917 15144 29929 15147
rect 29420 15116 29929 15144
rect 29420 15104 29426 15116
rect 29917 15113 29929 15116
rect 29963 15113 29975 15147
rect 29917 15107 29975 15113
rect 4341 15011 4399 15017
rect 4341 15008 4353 15011
rect 3436 14980 4353 15008
rect 3436 14949 3464 14980
rect 4341 14977 4353 14980
rect 4387 14977 4399 15011
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 4341 14971 4399 14977
rect 5828 14980 6745 15008
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2363 14912 2513 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14940 2651 14943
rect 2777 14943 2835 14949
rect 2777 14940 2789 14943
rect 2639 14912 2789 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 2777 14909 2789 14912
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 2915 14912 3341 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 3329 14909 3341 14912
rect 3375 14909 3387 14943
rect 3329 14903 3387 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3927 14912 4077 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 4154 14900 4160 14952
rect 4212 14900 4218 14952
rect 5828 14949 5856 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 7607 14980 7788 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14940 4491 14943
rect 4617 14943 4675 14949
rect 4617 14940 4629 14943
rect 4479 14912 4629 14940
rect 4479 14909 4491 14912
rect 4433 14903 4491 14909
rect 4617 14909 4629 14912
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14940 4767 14943
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4755 14912 4905 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5031 14912 5181 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5307 14912 5457 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5445 14909 5457 14912
rect 5491 14909 5503 14943
rect 5445 14903 5503 14909
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5583 14912 5733 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 5721 14909 5733 14912
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14909 5871 14943
rect 5813 14903 5871 14909
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6273 14943 6331 14949
rect 6273 14940 6285 14943
rect 6135 14912 6285 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6273 14909 6285 14912
rect 6319 14909 6331 14943
rect 6273 14903 6331 14909
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14940 6423 14943
rect 6454 14940 6460 14952
rect 6411 14912 6460 14940
rect 6411 14909 6423 14912
rect 6365 14903 6423 14909
rect 6454 14900 6460 14912
rect 6512 14900 6518 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 7101 14943 7159 14949
rect 7101 14940 7113 14943
rect 6871 14912 7113 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7101 14909 7113 14912
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 7208 14872 7236 14903
rect 7650 14900 7656 14952
rect 7708 14900 7714 14952
rect 7760 14949 7788 14980
rect 9232 14980 9413 15008
rect 9232 14949 9260 14980
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 9401 14971 9459 14977
rect 14752 14980 14933 15008
rect 7745 14943 7803 14949
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9306 14900 9312 14952
rect 9364 14900 9370 14952
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10468 14912 10701 14940
rect 10468 14900 10474 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 14752 14949 14780 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 14921 14971 14979 14977
rect 17144 14980 17325 15008
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11572 14912 11713 14940
rect 11572 14900 11578 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 14461 14943 14519 14949
rect 14461 14909 14473 14943
rect 14507 14940 14519 14943
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14507 14912 14657 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 17144 14949 17172 14980
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 18463 14980 18736 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 16577 14943 16635 14949
rect 16577 14909 16589 14943
rect 16623 14940 16635 14943
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16623 14912 16773 14940
rect 16623 14909 16635 14912
rect 16577 14903 16635 14909
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16761 14903 16819 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 16899 14912 17049 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17218 14900 17224 14952
rect 17276 14900 17282 14952
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 18598 14940 18604 14952
rect 18555 14912 18604 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18708 14949 18736 14980
rect 22664 14980 22845 15008
rect 22664 14949 22692 14980
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 23293 15011 23351 15017
rect 23293 14977 23305 15011
rect 23339 15008 23351 15011
rect 23339 14980 24348 15008
rect 23339 14977 23351 14980
rect 23293 14971 23351 14977
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 18785 14943 18843 14949
rect 18785 14909 18797 14943
rect 18831 14940 18843 14943
rect 18969 14943 19027 14949
rect 18969 14940 18981 14943
rect 18831 14912 18981 14940
rect 18831 14909 18843 14912
rect 18785 14903 18843 14909
rect 18969 14909 18981 14912
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14940 19119 14943
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 19107 14912 19257 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14940 19395 14943
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 19383 14912 19533 14940
rect 19383 14909 19395 14912
rect 19337 14903 19395 14909
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 19521 14903 19579 14909
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 20487 14912 20637 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 20625 14909 20637 14912
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 20717 14943 20775 14949
rect 20717 14909 20729 14943
rect 20763 14940 20775 14943
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20763 14912 20913 14940
rect 20763 14909 20775 14912
rect 20717 14903 20775 14909
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 20993 14943 21051 14949
rect 20993 14909 21005 14943
rect 21039 14940 21051 14943
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 21039 14912 21189 14940
rect 21039 14909 21051 14912
rect 20993 14903 21051 14909
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14940 21327 14943
rect 21453 14943 21511 14949
rect 21453 14940 21465 14943
rect 21315 14912 21465 14940
rect 21315 14909 21327 14912
rect 21269 14903 21327 14909
rect 21453 14909 21465 14912
rect 21499 14909 21511 14943
rect 21453 14903 21511 14909
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14940 21603 14943
rect 21729 14943 21787 14949
rect 21729 14940 21741 14943
rect 21591 14912 21741 14940
rect 21591 14909 21603 14912
rect 21545 14903 21603 14909
rect 21729 14909 21741 14912
rect 21775 14909 21787 14943
rect 21729 14903 21787 14909
rect 21821 14943 21879 14949
rect 21821 14909 21833 14943
rect 21867 14940 21879 14943
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 21867 14912 22017 14940
rect 21867 14909 21879 14912
rect 21821 14903 21879 14909
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22143 14912 22293 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 22373 14943 22431 14949
rect 22373 14909 22385 14943
rect 22419 14940 22431 14943
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 22419 14912 22569 14940
rect 22419 14909 22431 14912
rect 22373 14903 22431 14909
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 22738 14900 22744 14952
rect 22796 14900 22802 14952
rect 23385 14943 23443 14949
rect 23385 14909 23397 14943
rect 23431 14940 23443 14943
rect 23569 14943 23627 14949
rect 23569 14940 23581 14943
rect 23431 14912 23581 14940
rect 23431 14909 23443 14912
rect 23385 14903 23443 14909
rect 23569 14909 23581 14912
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 23658 14900 23664 14952
rect 23716 14900 23722 14952
rect 24320 14949 24348 14980
rect 24213 14943 24271 14949
rect 24213 14909 24225 14943
rect 24259 14909 24271 14943
rect 24213 14903 24271 14909
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24397 14943 24455 14949
rect 24397 14909 24409 14943
rect 24443 14940 24455 14943
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 24443 14912 24593 14940
rect 24443 14909 24455 14912
rect 24397 14903 24455 14909
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 7208 14844 7849 14872
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 24228 14872 24256 14903
rect 28994 14900 29000 14952
rect 29052 14900 29058 14952
rect 29089 14943 29147 14949
rect 29089 14909 29101 14943
rect 29135 14940 29147 14943
rect 29273 14943 29331 14949
rect 29273 14940 29285 14943
rect 29135 14912 29285 14940
rect 29135 14909 29147 14912
rect 29089 14903 29147 14909
rect 29273 14909 29285 14912
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 29365 14943 29423 14949
rect 29365 14909 29377 14943
rect 29411 14940 29423 14943
rect 29549 14943 29607 14949
rect 29549 14940 29561 14943
rect 29411 14912 29561 14940
rect 29411 14909 29423 14912
rect 29365 14903 29423 14909
rect 29549 14909 29561 14912
rect 29595 14909 29607 14943
rect 29549 14903 29607 14909
rect 29641 14943 29699 14949
rect 29641 14909 29653 14943
rect 29687 14940 29699 14943
rect 29825 14943 29883 14949
rect 29825 14940 29837 14943
rect 29687 14912 29837 14940
rect 29687 14909 29699 14912
rect 29641 14903 29699 14909
rect 29825 14909 29837 14912
rect 29871 14909 29883 14943
rect 29825 14903 29883 14909
rect 30561 14943 30619 14949
rect 30561 14909 30573 14943
rect 30607 14940 30619 14943
rect 31018 14940 31024 14952
rect 30607 14912 31024 14940
rect 30607 14909 30619 14912
rect 30561 14903 30619 14909
rect 31018 14900 31024 14912
rect 31076 14900 31082 14952
rect 24673 14875 24731 14881
rect 24673 14872 24685 14875
rect 24228 14844 24685 14872
rect 7837 14835 7895 14841
rect 24673 14841 24685 14844
rect 24719 14841 24731 14875
rect 24673 14835 24731 14841
rect 2225 14807 2283 14813
rect 2225 14773 2237 14807
rect 2271 14804 2283 14807
rect 2774 14804 2780 14816
rect 2271 14776 2780 14804
rect 2271 14773 2283 14776
rect 2225 14767 2283 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9214 14804 9220 14816
rect 9171 14776 9220 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 10870 14804 10876 14816
rect 10827 14776 10876 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 11388 14776 11805 14804
rect 11388 14764 11394 14776
rect 11793 14773 11805 14776
rect 11839 14773 11851 14807
rect 11793 14767 11851 14773
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16485 14807 16543 14813
rect 16485 14804 16497 14807
rect 16448 14776 16497 14804
rect 16448 14764 16454 14776
rect 16485 14773 16497 14776
rect 16531 14773 16543 14807
rect 16485 14767 16543 14773
rect 20349 14807 20407 14813
rect 20349 14773 20361 14807
rect 20395 14804 20407 14807
rect 20806 14804 20812 14816
rect 20395 14776 20812 14804
rect 20395 14773 20407 14776
rect 20349 14767 20407 14773
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 24118 14764 24124 14816
rect 24176 14764 24182 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 30469 14807 30527 14813
rect 30469 14804 30481 14807
rect 30432 14776 30481 14804
rect 30432 14764 30438 14776
rect 30469 14773 30481 14776
rect 30515 14773 30527 14807
rect 30469 14767 30527 14773
rect 552 14714 31648 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31648 14714
rect 552 14640 31648 14662
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 1872 14572 2881 14600
rect 1872 14473 1900 14572
rect 2869 14569 2881 14572
rect 2915 14569 2927 14603
rect 2869 14563 2927 14569
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4341 14603 4399 14609
rect 4341 14600 4353 14603
rect 4212 14572 4353 14600
rect 4212 14560 4218 14572
rect 4341 14569 4353 14572
rect 4387 14569 4399 14603
rect 4341 14563 4399 14569
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 7650 14560 7656 14612
rect 7708 14560 7714 14612
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 11514 14560 11520 14612
rect 11572 14560 11578 14612
rect 18598 14560 18604 14612
rect 18656 14560 18662 14612
rect 22094 14560 22100 14612
rect 22152 14560 22158 14612
rect 28994 14560 29000 14612
rect 29052 14600 29058 14612
rect 29089 14603 29147 14609
rect 29089 14600 29101 14603
rect 29052 14572 29101 14600
rect 29052 14560 29058 14572
rect 29089 14569 29101 14572
rect 29135 14569 29147 14603
rect 29089 14563 29147 14569
rect 31018 14560 31024 14612
rect 31076 14560 31082 14612
rect 2593 14535 2651 14541
rect 2593 14532 2605 14535
rect 2424 14504 2605 14532
rect 2424 14473 2452 14504
rect 2593 14501 2605 14504
rect 2639 14501 2651 14535
rect 2593 14495 2651 14501
rect 9033 14535 9091 14541
rect 9033 14501 9045 14535
rect 9079 14532 9091 14535
rect 14829 14535 14887 14541
rect 14829 14532 14841 14535
rect 9079 14504 9536 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2179 14436 2329 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14433 2467 14467
rect 2409 14427 2467 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 2516 14396 2544 14427
rect 2774 14424 2780 14476
rect 2832 14424 2838 14476
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 1811 14368 2544 14396
rect 4065 14399 4123 14405
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 4065 14365 4077 14399
rect 4111 14396 4123 14399
rect 4264 14396 4292 14427
rect 6086 14424 6092 14476
rect 6144 14424 6150 14476
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6365 14467 6423 14473
rect 6365 14464 6377 14467
rect 6227 14436 6377 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6365 14433 6377 14436
rect 6411 14433 6423 14467
rect 6365 14427 6423 14433
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14464 7803 14467
rect 7929 14467 7987 14473
rect 7929 14464 7941 14467
rect 7791 14436 7941 14464
rect 7791 14433 7803 14436
rect 7745 14427 7803 14433
rect 7929 14433 7941 14436
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14464 8079 14467
rect 8205 14467 8263 14473
rect 8205 14464 8217 14467
rect 8067 14436 8217 14464
rect 8067 14433 8079 14436
rect 8021 14427 8079 14433
rect 8205 14433 8217 14436
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14464 8355 14467
rect 8481 14467 8539 14473
rect 8481 14464 8493 14467
rect 8343 14436 8493 14464
rect 8343 14433 8355 14436
rect 8297 14427 8355 14433
rect 8481 14433 8493 14436
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 8619 14436 8769 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 8849 14467 8907 14473
rect 8849 14433 8861 14467
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 4111 14368 4292 14396
rect 4111 14365 4123 14368
rect 4065 14359 4123 14365
rect 8864 14328 8892 14427
rect 9140 14396 9168 14427
rect 9214 14424 9220 14476
rect 9272 14424 9278 14476
rect 9508 14473 9536 14504
rect 14108 14504 14841 14532
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10689 14467 10747 14473
rect 10689 14464 10701 14467
rect 10551 14436 10701 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10689 14433 10701 14436
rect 10735 14433 10747 14467
rect 10689 14427 10747 14433
rect 10778 14424 10784 14476
rect 10836 14424 10842 14476
rect 11330 14424 11336 14476
rect 11388 14424 11394 14476
rect 14108 14473 14136 14504
rect 14829 14501 14841 14504
rect 14875 14501 14887 14535
rect 14829 14495 14887 14501
rect 16301 14535 16359 14541
rect 16301 14501 16313 14535
rect 16347 14532 16359 14535
rect 22925 14535 22983 14541
rect 22925 14532 22937 14535
rect 16347 14504 16528 14532
rect 16347 14501 16359 14504
rect 16301 14495 16359 14501
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11655 14436 11805 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11931 14436 12081 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12161 14467 12219 14473
rect 12161 14433 12173 14467
rect 12207 14464 12219 14467
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12207 14436 12357 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12621 14467 12679 14473
rect 12621 14464 12633 14467
rect 12483 14436 12633 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12621 14433 12633 14436
rect 12667 14433 12679 14467
rect 12621 14427 12679 14433
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 12897 14467 12955 14473
rect 12897 14464 12909 14467
rect 12759 14436 12909 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 12897 14433 12909 14436
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 13035 14436 13185 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 13265 14467 13323 14473
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13449 14467 13507 14473
rect 13449 14464 13461 14467
rect 13311 14436 13461 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13449 14433 13461 14436
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13587 14436 13737 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 13725 14427 13783 14433
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13863 14436 14013 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 14001 14427 14059 14433
rect 14093 14467 14151 14473
rect 14093 14433 14105 14467
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14366 14424 14372 14476
rect 14424 14424 14430 14476
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14599 14436 14749 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 14737 14433 14749 14436
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15427 14436 15577 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14464 15715 14467
rect 15841 14467 15899 14473
rect 15841 14464 15853 14467
rect 15703 14436 15853 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 15841 14433 15853 14436
rect 15887 14433 15899 14467
rect 15841 14427 15899 14433
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 9140 14368 9321 14396
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 14476 14396 14504 14427
rect 14323 14368 14504 14396
rect 15948 14396 15976 14427
rect 16390 14424 16396 14476
rect 16448 14424 16454 14476
rect 16500 14473 16528 14504
rect 22204 14504 22937 14532
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 17586 14424 17592 14476
rect 17644 14424 17650 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 17773 14467 17831 14473
rect 17773 14433 17785 14467
rect 17819 14464 17831 14467
rect 17957 14467 18015 14473
rect 17957 14464 17969 14467
rect 17819 14436 17969 14464
rect 17819 14433 17831 14436
rect 17773 14427 17831 14433
rect 17957 14433 17969 14436
rect 18003 14433 18015 14467
rect 17957 14427 18015 14433
rect 18049 14467 18107 14473
rect 18049 14433 18061 14467
rect 18095 14464 18107 14467
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18095 14436 18245 14464
rect 18095 14433 18107 14436
rect 18049 14427 18107 14433
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14464 18383 14467
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 18371 14436 18521 14464
rect 18371 14433 18383 14436
rect 18325 14427 18383 14433
rect 18509 14433 18521 14436
rect 18555 14433 18567 14467
rect 18509 14427 18567 14433
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14464 20499 14467
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 20487 14436 20637 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 15948 14368 16589 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 16577 14365 16589 14368
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 17696 14396 17724 14427
rect 17543 14368 17724 14396
rect 20732 14396 20760 14427
rect 20806 14424 20812 14476
rect 20864 14424 20870 14476
rect 22204 14473 22232 14504
rect 22925 14501 22937 14504
rect 22971 14501 22983 14535
rect 22925 14495 22983 14501
rect 22189 14467 22247 14473
rect 22189 14433 22201 14467
rect 22235 14433 22247 14467
rect 22189 14427 22247 14433
rect 22462 14424 22468 14476
rect 22520 14424 22526 14476
rect 22557 14467 22615 14473
rect 22557 14433 22569 14467
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 22649 14467 22707 14473
rect 22649 14433 22661 14467
rect 22695 14464 22707 14467
rect 22833 14467 22891 14473
rect 22833 14464 22845 14467
rect 22695 14436 22845 14464
rect 22695 14433 22707 14436
rect 22649 14427 22707 14433
rect 22833 14433 22845 14436
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20732 14368 20913 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14396 22431 14399
rect 22572 14396 22600 14427
rect 24118 14424 24124 14476
rect 24176 14424 24182 14476
rect 24213 14467 24271 14473
rect 24213 14433 24225 14467
rect 24259 14433 24271 14467
rect 24213 14427 24271 14433
rect 24305 14467 24363 14473
rect 24305 14433 24317 14467
rect 24351 14464 24363 14467
rect 24489 14467 24547 14473
rect 24489 14464 24501 14467
rect 24351 14436 24501 14464
rect 24351 14433 24363 14436
rect 24305 14427 24363 14433
rect 24489 14433 24501 14436
rect 24535 14433 24547 14467
rect 24489 14427 24547 14433
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24765 14467 24823 14473
rect 24765 14464 24777 14467
rect 24627 14436 24777 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24765 14433 24777 14436
rect 24811 14433 24823 14467
rect 24765 14427 24823 14433
rect 24857 14467 24915 14473
rect 24857 14433 24869 14467
rect 24903 14464 24915 14467
rect 25041 14467 25099 14473
rect 25041 14464 25053 14467
rect 24903 14436 25053 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 25041 14433 25053 14436
rect 25087 14433 25099 14467
rect 25041 14427 25099 14433
rect 29181 14467 29239 14473
rect 29181 14433 29193 14467
rect 29227 14464 29239 14467
rect 29365 14467 29423 14473
rect 29365 14464 29377 14467
rect 29227 14436 29377 14464
rect 29227 14433 29239 14436
rect 29181 14427 29239 14433
rect 29365 14433 29377 14436
rect 29411 14433 29423 14467
rect 29365 14427 29423 14433
rect 29457 14467 29515 14473
rect 29457 14433 29469 14467
rect 29503 14464 29515 14467
rect 29641 14467 29699 14473
rect 29641 14464 29653 14467
rect 29503 14436 29653 14464
rect 29503 14433 29515 14436
rect 29457 14427 29515 14433
rect 29641 14433 29653 14436
rect 29687 14433 29699 14467
rect 29641 14427 29699 14433
rect 29733 14467 29791 14473
rect 29733 14433 29745 14467
rect 29779 14464 29791 14467
rect 29917 14467 29975 14473
rect 29917 14464 29929 14467
rect 29779 14436 29929 14464
rect 29779 14433 29791 14436
rect 29733 14427 29791 14433
rect 29917 14433 29929 14436
rect 29963 14433 29975 14467
rect 29917 14427 29975 14433
rect 30009 14467 30067 14473
rect 30009 14433 30021 14467
rect 30055 14464 30067 14467
rect 30193 14467 30251 14473
rect 30193 14464 30205 14467
rect 30055 14436 30205 14464
rect 30055 14433 30067 14436
rect 30009 14427 30067 14433
rect 30193 14433 30205 14436
rect 30239 14433 30251 14467
rect 30193 14427 30251 14433
rect 30285 14467 30343 14473
rect 30285 14433 30297 14467
rect 30331 14433 30343 14467
rect 30285 14427 30343 14433
rect 22419 14368 22600 14396
rect 24029 14399 24087 14405
rect 22419 14365 22431 14368
rect 22373 14359 22431 14365
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 24228 14396 24256 14427
rect 24075 14368 24256 14396
rect 30300 14396 30328 14427
rect 30374 14424 30380 14476
rect 30432 14424 30438 14476
rect 30834 14424 30840 14476
rect 30892 14424 30898 14476
rect 30929 14467 30987 14473
rect 30929 14433 30941 14467
rect 30975 14433 30987 14467
rect 30929 14427 30987 14433
rect 30469 14399 30527 14405
rect 30469 14396 30481 14399
rect 30300 14368 30481 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 30469 14365 30481 14368
rect 30515 14365 30527 14399
rect 30469 14359 30527 14365
rect 30745 14399 30803 14405
rect 30745 14365 30757 14399
rect 30791 14396 30803 14399
rect 30944 14396 30972 14427
rect 30791 14368 30972 14396
rect 30791 14365 30803 14368
rect 30745 14359 30803 14365
rect 9585 14331 9643 14337
rect 9585 14328 9597 14331
rect 8864 14300 9597 14328
rect 9585 14297 9597 14300
rect 9631 14297 9643 14331
rect 9585 14291 9643 14297
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14260 2099 14263
rect 2498 14260 2504 14272
rect 2087 14232 2504 14260
rect 2087 14229 2099 14232
rect 2041 14223 2099 14229
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 16206 14260 16212 14272
rect 15335 14232 16212 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 20349 14263 20407 14269
rect 20349 14260 20361 14263
rect 20312 14232 20361 14260
rect 20312 14220 20318 14232
rect 20349 14229 20361 14232
rect 20395 14229 20407 14263
rect 20349 14223 20407 14229
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 552 14170 31648 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31648 14170
rect 552 14096 31648 14118
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4212 14028 4905 14056
rect 4212 14016 4218 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 4893 14019 4951 14025
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10836 14028 11345 14056
rect 10836 14016 10842 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17644 14028 17785 14056
rect 17644 14016 17650 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 23201 14059 23259 14065
rect 23201 14056 23213 14059
rect 22520 14028 23213 14056
rect 22520 14016 22526 14028
rect 23201 14025 23213 14028
rect 23247 14025 23259 14059
rect 23201 14019 23259 14025
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 31113 14059 31171 14065
rect 31113 14056 31125 14059
rect 30892 14028 31125 14056
rect 30892 14016 30898 14028
rect 31113 14025 31125 14028
rect 31159 14025 31171 14059
rect 31113 14019 31171 14025
rect 19153 13991 19211 13997
rect 19153 13957 19165 13991
rect 19199 13988 19211 13991
rect 19426 13988 19432 14000
rect 19199 13960 19432 13988
rect 19199 13957 19211 13960
rect 19153 13951 19211 13957
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2424 13892 2605 13920
rect 2424 13861 2452 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 2593 13883 2651 13889
rect 6472 13892 7021 13920
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 2179 13824 2329 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 2498 13812 2504 13864
rect 2556 13812 2562 13864
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 6472 13861 6500 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 16301 13923 16359 13929
rect 16301 13920 16313 13923
rect 7009 13883 7067 13889
rect 16132 13892 16313 13920
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 4111 13824 4261 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4387 13824 4537 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4663 13824 4813 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5951 13824 6101 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6227 13824 6377 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6365 13815 6423 13821
rect 6457 13855 6515 13861
rect 6457 13821 6469 13855
rect 6503 13821 6515 13855
rect 6457 13815 6515 13821
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6779 13824 6929 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10643 13824 10793 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 10870 13812 10876 13864
rect 10928 13812 10934 13864
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 16132 13861 16160 13892
rect 16301 13889 16313 13892
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13920 17279 13923
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 17267 13892 17448 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 15749 13855 15807 13861
rect 15749 13852 15761 13855
rect 15611 13824 15761 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 15749 13821 15761 13824
rect 15795 13821 15807 13855
rect 15749 13815 15807 13821
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15887 13824 16037 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16025 13821 16037 13824
rect 16071 13821 16083 13855
rect 16025 13815 16083 13821
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 17310 13812 17316 13864
rect 17368 13812 17374 13864
rect 17420 13861 17448 13892
rect 20916 13892 21097 13920
rect 20916 13861 20944 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 25041 13923 25099 13929
rect 22143 13892 22324 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 17681 13855 17739 13861
rect 17681 13852 17693 13855
rect 17543 13824 17693 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 17681 13821 17693 13824
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19429 13855 19487 13861
rect 19429 13852 19441 13855
rect 19291 13824 19441 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19429 13821 19441 13824
rect 19475 13821 19487 13855
rect 19429 13815 19487 13821
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13852 19579 13855
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19567 13824 19717 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13852 19855 13855
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19843 13824 19993 13852
rect 19843 13821 19855 13824
rect 19797 13815 19855 13821
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20257 13855 20315 13861
rect 20257 13852 20269 13855
rect 20119 13824 20269 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20257 13821 20269 13824
rect 20303 13821 20315 13855
rect 20257 13815 20315 13821
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20395 13824 20545 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20671 13824 20821 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 22186 13812 22192 13864
rect 22244 13812 22250 13864
rect 22296 13861 22324 13892
rect 25041 13889 25053 13923
rect 25087 13920 25099 13923
rect 30561 13923 30619 13929
rect 25087 13892 25268 13920
rect 25087 13889 25099 13892
rect 25041 13883 25099 13889
rect 22281 13855 22339 13861
rect 22281 13821 22293 13855
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 22419 13824 22569 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 22557 13821 22569 13824
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22695 13824 22845 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 22925 13855 22983 13861
rect 22925 13821 22937 13855
rect 22971 13852 22983 13855
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 22971 13824 23121 13852
rect 22971 13821 22983 13824
rect 22925 13815 22983 13821
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 25130 13812 25136 13864
rect 25188 13812 25194 13864
rect 25240 13861 25268 13892
rect 30561 13889 30573 13923
rect 30607 13920 30619 13923
rect 30607 13892 30788 13920
rect 30607 13889 30619 13892
rect 30561 13883 30619 13889
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 25317 13855 25375 13861
rect 25317 13821 25329 13855
rect 25363 13852 25375 13855
rect 25501 13855 25559 13861
rect 25501 13852 25513 13855
rect 25363 13824 25513 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 25501 13821 25513 13824
rect 25547 13821 25559 13855
rect 25501 13815 25559 13821
rect 25593 13855 25651 13861
rect 25593 13821 25605 13855
rect 25639 13852 25651 13855
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25639 13824 25789 13852
rect 25639 13821 25651 13824
rect 25593 13815 25651 13821
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 26053 13855 26111 13861
rect 26053 13852 26065 13855
rect 25915 13824 26065 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 26053 13821 26065 13824
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 26329 13855 26387 13861
rect 26329 13852 26341 13855
rect 26191 13824 26341 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 26329 13821 26341 13824
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 26421 13855 26479 13861
rect 26421 13821 26433 13855
rect 26467 13852 26479 13855
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 26467 13824 26617 13852
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 26605 13821 26617 13824
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 26697 13855 26755 13861
rect 26697 13821 26709 13855
rect 26743 13852 26755 13855
rect 26881 13855 26939 13861
rect 26881 13852 26893 13855
rect 26743 13824 26893 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 26881 13821 26893 13824
rect 26927 13821 26939 13855
rect 26881 13815 26939 13821
rect 26973 13855 27031 13861
rect 26973 13821 26985 13855
rect 27019 13852 27031 13855
rect 27157 13855 27215 13861
rect 27157 13852 27169 13855
rect 27019 13824 27169 13852
rect 27019 13821 27031 13824
rect 26973 13815 27031 13821
rect 27157 13821 27169 13824
rect 27203 13821 27215 13855
rect 27157 13815 27215 13821
rect 27249 13855 27307 13861
rect 27249 13821 27261 13855
rect 27295 13852 27307 13855
rect 27433 13855 27491 13861
rect 27433 13852 27445 13855
rect 27295 13824 27445 13852
rect 27295 13821 27307 13824
rect 27249 13815 27307 13821
rect 27433 13821 27445 13824
rect 27479 13821 27491 13855
rect 27433 13815 27491 13821
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13852 27583 13855
rect 27709 13855 27767 13861
rect 27709 13852 27721 13855
rect 27571 13824 27721 13852
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 27709 13821 27721 13824
rect 27755 13821 27767 13855
rect 27709 13815 27767 13821
rect 27801 13855 27859 13861
rect 27801 13821 27813 13855
rect 27847 13852 27859 13855
rect 27985 13855 28043 13861
rect 27985 13852 27997 13855
rect 27847 13824 27997 13852
rect 27847 13821 27859 13824
rect 27801 13815 27859 13821
rect 27985 13821 27997 13824
rect 28031 13821 28043 13855
rect 27985 13815 28043 13821
rect 28077 13855 28135 13861
rect 28077 13821 28089 13855
rect 28123 13852 28135 13855
rect 28261 13855 28319 13861
rect 28261 13852 28273 13855
rect 28123 13824 28273 13852
rect 28123 13821 28135 13824
rect 28077 13815 28135 13821
rect 28261 13821 28273 13824
rect 28307 13821 28319 13855
rect 28261 13815 28319 13821
rect 28353 13855 28411 13861
rect 28353 13821 28365 13855
rect 28399 13852 28411 13855
rect 28537 13855 28595 13861
rect 28537 13852 28549 13855
rect 28399 13824 28549 13852
rect 28399 13821 28411 13824
rect 28353 13815 28411 13821
rect 28537 13821 28549 13824
rect 28583 13821 28595 13855
rect 28537 13815 28595 13821
rect 28629 13855 28687 13861
rect 28629 13821 28641 13855
rect 28675 13852 28687 13855
rect 28997 13855 29055 13861
rect 28997 13852 29009 13855
rect 28675 13824 29009 13852
rect 28675 13821 28687 13824
rect 28629 13815 28687 13821
rect 28997 13821 29009 13824
rect 29043 13821 29055 13855
rect 28997 13815 29055 13821
rect 30650 13812 30656 13864
rect 30708 13812 30714 13864
rect 30760 13861 30788 13892
rect 30745 13855 30803 13861
rect 30745 13821 30757 13855
rect 30791 13821 30803 13855
rect 30745 13815 30803 13821
rect 30837 13855 30895 13861
rect 30837 13821 30849 13855
rect 30883 13852 30895 13855
rect 31021 13855 31079 13861
rect 31021 13852 31033 13855
rect 30883 13824 31033 13852
rect 30883 13821 30895 13824
rect 30837 13815 30895 13821
rect 31021 13821 31033 13824
rect 31067 13821 31079 13855
rect 31021 13815 31079 13821
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2041 13719 2099 13725
rect 2041 13716 2053 13719
rect 2004 13688 2053 13716
rect 2004 13676 2010 13688
rect 2041 13685 2053 13688
rect 2087 13685 2099 13719
rect 2041 13679 2099 13685
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 6086 13716 6092 13728
rect 5859 13688 6092 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10962 13716 10968 13728
rect 10551 13688 10968 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11664 13688 11897 13716
rect 11664 13676 11670 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 11885 13679 11943 13685
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15473 13719 15531 13725
rect 15473 13716 15485 13719
rect 15344 13688 15485 13716
rect 15344 13676 15350 13688
rect 15473 13685 15485 13688
rect 15519 13685 15531 13719
rect 15473 13679 15531 13685
rect 29086 13676 29092 13728
rect 29144 13676 29150 13728
rect 552 13626 31648 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31648 13626
rect 552 13552 31648 13574
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 4028 13484 4077 13512
rect 4028 13472 4034 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 6178 13472 6184 13524
rect 6236 13472 6242 13524
rect 6638 13472 6644 13524
rect 6696 13472 6702 13524
rect 11790 13472 11796 13524
rect 11848 13472 11854 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17368 13484 17877 13512
rect 17368 13472 17374 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 20349 13515 20407 13521
rect 20349 13481 20361 13515
rect 20395 13512 20407 13515
rect 20990 13512 20996 13524
rect 20395 13484 20996 13512
rect 20395 13481 20407 13484
rect 20349 13475 20407 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22741 13515 22799 13521
rect 22741 13512 22753 13515
rect 22244 13484 22753 13512
rect 22244 13472 22250 13484
rect 22741 13481 22753 13484
rect 22787 13481 22799 13515
rect 22741 13475 22799 13481
rect 30650 13472 30656 13524
rect 30708 13512 30714 13524
rect 31205 13515 31263 13521
rect 31205 13512 31217 13515
rect 30708 13484 31217 13512
rect 30708 13472 30714 13484
rect 31205 13481 31217 13484
rect 31251 13481 31263 13515
rect 31205 13475 31263 13481
rect 1857 13447 1915 13453
rect 1857 13413 1869 13447
rect 1903 13444 1915 13447
rect 2961 13447 3019 13453
rect 2961 13444 2973 13447
rect 1903 13416 2084 13444
rect 1903 13413 1915 13416
rect 1857 13407 1915 13413
rect 1946 13336 1952 13388
rect 2004 13336 2010 13388
rect 2056 13385 2084 13416
rect 2792 13416 2973 13444
rect 2792 13385 2820 13416
rect 2961 13413 2973 13416
rect 3007 13413 3019 13447
rect 4893 13447 4951 13453
rect 4893 13444 4905 13447
rect 2961 13407 3019 13413
rect 4172 13416 4905 13444
rect 4172 13385 4200 13416
rect 4893 13413 4905 13416
rect 4939 13413 4951 13447
rect 4893 13407 4951 13413
rect 12989 13447 13047 13453
rect 12989 13413 13001 13447
rect 13035 13444 13047 13447
rect 15197 13447 15255 13453
rect 13035 13416 13216 13444
rect 13035 13413 13047 13416
rect 12989 13407 13047 13413
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2547 13348 2697 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2884 13308 2912 13339
rect 4246 13336 4252 13388
rect 4304 13336 4310 13388
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4387 13348 4537 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4663 13348 4813 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 6086 13336 6092 13388
rect 6144 13336 6150 13388
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6779 13348 6929 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 7006 13336 7012 13388
rect 7064 13336 7070 13388
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7331 13348 7481 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 7607 13348 7757 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 7745 13345 7757 13348
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13376 7895 13379
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7883 13348 8033 13376
rect 7883 13345 7895 13348
rect 7837 13339 7895 13345
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 8159 13348 8309 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 8435 13348 8585 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8573 13345 8585 13348
rect 8619 13345 8631 13379
rect 8573 13339 8631 13345
rect 8665 13379 8723 13385
rect 8665 13345 8677 13379
rect 8711 13376 8723 13379
rect 8849 13379 8907 13385
rect 8849 13376 8861 13379
rect 8711 13348 8861 13376
rect 8711 13345 8723 13348
rect 8665 13339 8723 13345
rect 8849 13345 8861 13348
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8987 13348 9137 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9263 13348 9413 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9539 13348 9689 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9815 13348 9965 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10091 13348 10241 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10367 13348 10517 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 2179 13280 2912 13308
rect 10612 13308 10640 13339
rect 10962 13336 10968 13388
rect 11020 13336 11026 13388
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13376 11943 13379
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11931 13348 12081 13376
rect 11931 13345 11943 13348
rect 11885 13339 11943 13345
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13376 12219 13379
rect 12345 13379 12403 13385
rect 12345 13376 12357 13379
rect 12207 13348 12357 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 12345 13345 12357 13348
rect 12391 13345 12403 13379
rect 12345 13339 12403 13345
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12483 13348 12633 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 11057 13311 11115 13317
rect 11057 13308 11069 13311
rect 10612 13280 11069 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 11057 13277 11069 13280
rect 11103 13277 11115 13311
rect 12728 13308 12756 13339
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 13188 13385 13216 13416
rect 15197 13413 15209 13447
rect 15243 13444 15255 13447
rect 18141 13447 18199 13453
rect 18141 13444 18153 13447
rect 15243 13416 16160 13444
rect 15243 13413 15255 13416
rect 15197 13407 15255 13413
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 15286 13336 15292 13388
rect 15344 13336 15350 13388
rect 16132 13385 16160 13416
rect 17420 13416 18153 13444
rect 17420 13385 17448 13416
rect 18141 13413 18153 13416
rect 18187 13413 18199 13447
rect 18141 13407 18199 13413
rect 15565 13379 15623 13385
rect 15565 13345 15577 13379
rect 15611 13376 15623 13379
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15611 13348 15761 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13345 17463 13379
rect 17405 13339 17463 13345
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13376 17647 13379
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 17635 13348 17785 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 18233 13379 18291 13385
rect 18233 13345 18245 13379
rect 18279 13376 18291 13379
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 18279 13348 18429 13376
rect 18279 13345 18291 13348
rect 18233 13339 18291 13345
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 18417 13339 18475 13345
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18555 13348 18705 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13376 18843 13379
rect 18969 13379 19027 13385
rect 18969 13376 18981 13379
rect 18831 13348 18981 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 18969 13345 18981 13348
rect 19015 13345 19027 13379
rect 18969 13339 19027 13345
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13376 19119 13379
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 19107 13348 19257 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13345 19395 13379
rect 19337 13339 19395 13345
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 12728 13280 13277 13308
rect 11057 13271 11115 13277
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 15856 13308 15884 13339
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15856 13280 16221 13308
rect 13265 13271 13323 13277
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17512 13308 17540 13339
rect 17359 13280 17540 13308
rect 19352 13308 19380 13339
rect 19426 13336 19432 13388
rect 19484 13336 19490 13388
rect 20254 13336 20260 13388
rect 20312 13336 20318 13388
rect 21542 13336 21548 13388
rect 21600 13336 21606 13388
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13376 21695 13379
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21683 13348 21833 13376
rect 21683 13345 21695 13348
rect 21637 13339 21695 13345
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 21913 13379 21971 13385
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22097 13379 22155 13385
rect 22097 13376 22109 13379
rect 21959 13348 22109 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22097 13345 22109 13348
rect 22143 13345 22155 13379
rect 22097 13339 22155 13345
rect 22189 13379 22247 13385
rect 22189 13345 22201 13379
rect 22235 13376 22247 13379
rect 22373 13379 22431 13385
rect 22373 13376 22385 13379
rect 22235 13348 22385 13376
rect 22235 13345 22247 13348
rect 22189 13339 22247 13345
rect 22373 13345 22385 13348
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 22465 13379 22523 13385
rect 22465 13345 22477 13379
rect 22511 13376 22523 13379
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22511 13348 22661 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25087 13348 25237 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 25225 13345 25237 13348
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13376 25375 13379
rect 25593 13379 25651 13385
rect 25593 13376 25605 13379
rect 25363 13348 25605 13376
rect 25363 13345 25375 13348
rect 25317 13339 25375 13345
rect 25593 13345 25605 13348
rect 25639 13345 25651 13379
rect 25593 13339 25651 13345
rect 25685 13379 25743 13385
rect 25685 13345 25697 13379
rect 25731 13376 25743 13379
rect 25869 13379 25927 13385
rect 25869 13376 25881 13379
rect 25731 13348 25881 13376
rect 25731 13345 25743 13348
rect 25685 13339 25743 13345
rect 25869 13345 25881 13348
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 25961 13379 26019 13385
rect 25961 13345 25973 13379
rect 26007 13376 26019 13379
rect 26142 13376 26148 13388
rect 26007 13348 26148 13376
rect 26007 13345 26019 13348
rect 25961 13339 26019 13345
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 26602 13336 26608 13388
rect 26660 13336 26666 13388
rect 28445 13379 28503 13385
rect 28445 13345 28457 13379
rect 28491 13376 28503 13379
rect 28629 13379 28687 13385
rect 28629 13376 28641 13379
rect 28491 13348 28641 13376
rect 28491 13345 28503 13348
rect 28445 13339 28503 13345
rect 28629 13345 28641 13348
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 28721 13379 28779 13385
rect 28721 13345 28733 13379
rect 28767 13376 28779 13379
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 28767 13348 28917 13376
rect 28767 13345 28779 13348
rect 28721 13339 28779 13345
rect 28905 13345 28917 13348
rect 28951 13345 28963 13379
rect 28905 13339 28963 13345
rect 28997 13379 29055 13385
rect 28997 13345 29009 13379
rect 29043 13345 29055 13379
rect 28997 13339 29055 13345
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 19352 13280 19533 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 29012 13308 29040 13339
rect 29086 13336 29092 13388
rect 29144 13336 29150 13388
rect 30190 13336 30196 13388
rect 30248 13336 30254 13388
rect 30285 13379 30343 13385
rect 30285 13345 30297 13379
rect 30331 13345 30343 13379
rect 30285 13339 30343 13345
rect 30377 13379 30435 13385
rect 30377 13345 30389 13379
rect 30423 13376 30435 13379
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 30423 13348 30573 13376
rect 30423 13345 30435 13348
rect 30377 13339 30435 13345
rect 30561 13345 30573 13348
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 30653 13379 30711 13385
rect 30653 13345 30665 13379
rect 30699 13376 30711 13379
rect 30837 13379 30895 13385
rect 30837 13376 30849 13379
rect 30699 13348 30849 13376
rect 30699 13345 30711 13348
rect 30653 13339 30711 13345
rect 30837 13345 30849 13348
rect 30883 13345 30895 13379
rect 30837 13339 30895 13345
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13376 30987 13379
rect 31113 13379 31171 13385
rect 31113 13376 31125 13379
rect 30975 13348 31125 13376
rect 30975 13345 30987 13348
rect 30929 13339 30987 13345
rect 31113 13345 31125 13348
rect 31159 13345 31171 13379
rect 31113 13339 31171 13345
rect 29181 13311 29239 13317
rect 29181 13308 29193 13311
rect 29012 13280 29193 13308
rect 19521 13271 19579 13277
rect 29181 13277 29193 13280
rect 29227 13277 29239 13311
rect 29181 13271 29239 13277
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30300 13308 30328 13339
rect 30147 13280 30328 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 2406 13132 2412 13184
rect 2464 13132 2470 13184
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7374 13172 7380 13184
rect 7239 13144 7380 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 11974 13172 11980 13184
rect 11563 13144 11980 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 15654 13172 15660 13184
rect 15519 13144 15660 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 24949 13175 25007 13181
rect 24949 13141 24961 13175
rect 24995 13172 25007 13175
rect 25314 13172 25320 13184
rect 24995 13144 25320 13172
rect 24995 13141 25007 13144
rect 24949 13135 25007 13141
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 26513 13175 26571 13181
rect 26513 13141 26525 13175
rect 26559 13172 26571 13175
rect 26878 13172 26884 13184
rect 26559 13144 26884 13172
rect 26559 13141 26571 13144
rect 26513 13135 26571 13141
rect 26878 13132 26884 13144
rect 26936 13132 26942 13184
rect 28353 13175 28411 13181
rect 28353 13141 28365 13175
rect 28399 13172 28411 13175
rect 28994 13172 29000 13184
rect 28399 13144 29000 13172
rect 28399 13141 28411 13144
rect 28353 13135 28411 13141
rect 28994 13132 29000 13144
rect 29052 13132 29058 13184
rect 552 13082 31648 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31648 13082
rect 552 13008 31648 13030
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4246 12968 4252 12980
rect 4203 12940 4252 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 7064 12940 7481 12968
rect 7064 12928 7070 12940
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 7469 12931 7527 12937
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13136 12940 13921 12968
rect 13136 12928 13142 12940
rect 13909 12937 13921 12940
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 21542 12928 21548 12980
rect 21600 12968 21606 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 21600 12940 21649 12968
rect 21600 12928 21606 12940
rect 21637 12937 21649 12940
rect 21683 12937 21695 12971
rect 21637 12931 21695 12937
rect 26142 12928 26148 12980
rect 26200 12928 26206 12980
rect 26602 12928 26608 12980
rect 26660 12968 26666 12980
rect 26881 12971 26939 12977
rect 26881 12968 26893 12971
rect 26660 12940 26893 12968
rect 26660 12928 26666 12940
rect 26881 12937 26893 12940
rect 26927 12937 26939 12971
rect 26881 12931 26939 12937
rect 30190 12928 30196 12980
rect 30248 12968 30254 12980
rect 30745 12971 30803 12977
rect 30745 12968 30757 12971
rect 30248 12940 30757 12968
rect 30248 12928 30254 12940
rect 30745 12937 30757 12940
rect 30791 12937 30803 12971
rect 30745 12931 30803 12937
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2363 12804 2544 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2406 12724 2412 12776
rect 2464 12724 2470 12776
rect 2516 12773 2544 12804
rect 2976 12804 3341 12832
rect 2976 12773 3004 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 3329 12795 3387 12801
rect 4816 12804 5365 12832
rect 4816 12773 4844 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 13311 12804 13584 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12733 3019 12767
rect 2961 12727 3019 12733
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4295 12736 4445 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4571 12736 4721 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 2593 12699 2651 12705
rect 2593 12665 2605 12699
rect 2639 12696 2651 12699
rect 3252 12696 3280 12727
rect 4982 12724 4988 12776
rect 5040 12724 5046 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 5123 12736 5273 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12764 6239 12767
rect 6270 12764 6276 12776
rect 6227 12736 6276 12764
rect 6227 12733 6239 12736
rect 6181 12727 6239 12733
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 7374 12724 7380 12776
rect 7432 12724 7438 12776
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11655 12736 11805 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 11885 12767 11943 12773
rect 11885 12733 11897 12767
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 2639 12668 3280 12696
rect 11900 12696 11928 12727
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 13556 12773 13584 12804
rect 15580 12804 15761 12832
rect 15580 12773 15608 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 19107 12804 19288 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13679 12736 13829 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15335 12736 15485 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11900 12668 12081 12696
rect 2639 12665 2651 12668
rect 2593 12659 2651 12665
rect 12069 12665 12081 12668
rect 12115 12665 12127 12699
rect 13372 12696 13400 12727
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 19260 12773 19288 12804
rect 21744 12804 22477 12832
rect 21744 12773 21772 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 22465 12795 22523 12801
rect 25240 12804 25421 12832
rect 19153 12767 19211 12773
rect 19153 12733 19165 12767
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 19383 12736 19533 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19659 12736 19809 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 19797 12733 19809 12736
rect 19843 12733 19855 12767
rect 19797 12727 19855 12733
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19935 12736 20085 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 20165 12767 20223 12773
rect 20165 12733 20177 12767
rect 20211 12764 20223 12767
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 20211 12736 20361 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 21729 12767 21787 12773
rect 21729 12733 21741 12767
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 13906 12696 13912 12708
rect 13372 12668 13912 12696
rect 12069 12659 12127 12665
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 19168 12696 19196 12727
rect 21818 12724 21824 12776
rect 21876 12724 21882 12776
rect 25240 12773 25268 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 30834 12832 30840 12844
rect 26651 12804 26832 12832
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 21913 12767 21971 12773
rect 21913 12733 21925 12767
rect 21959 12764 21971 12767
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21959 12736 22109 12764
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12764 22247 12767
rect 22373 12767 22431 12773
rect 22373 12764 22385 12767
rect 22235 12736 22385 12764
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 22373 12733 22385 12736
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 24397 12767 24455 12773
rect 24397 12733 24409 12767
rect 24443 12764 24455 12767
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 24443 12736 24593 12764
rect 24443 12733 24455 12736
rect 24397 12727 24455 12733
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12764 24731 12767
rect 24857 12767 24915 12773
rect 24857 12764 24869 12767
rect 24719 12736 24869 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 24857 12733 24869 12736
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12764 25007 12767
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24995 12736 25145 12764
rect 24995 12733 25007 12736
rect 24949 12727 25007 12733
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12733 25283 12767
rect 25225 12727 25283 12733
rect 25314 12724 25320 12776
rect 25372 12724 25378 12776
rect 26237 12767 26295 12773
rect 26237 12733 26249 12767
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 19426 12696 19432 12708
rect 19168 12668 19432 12696
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 26252 12696 26280 12727
rect 26694 12724 26700 12776
rect 26752 12724 26758 12776
rect 26804 12773 26832 12804
rect 30024 12804 30840 12832
rect 26789 12767 26847 12773
rect 26789 12733 26801 12767
rect 26835 12733 26847 12767
rect 26789 12727 26847 12733
rect 26878 12724 26884 12776
rect 26936 12764 26942 12776
rect 27065 12767 27123 12773
rect 27065 12764 27077 12767
rect 26936 12736 27077 12764
rect 26936 12724 26942 12736
rect 27065 12733 27077 12736
rect 27111 12733 27123 12767
rect 27065 12727 27123 12733
rect 28353 12767 28411 12773
rect 28353 12733 28365 12767
rect 28399 12764 28411 12767
rect 28537 12767 28595 12773
rect 28537 12764 28549 12767
rect 28399 12736 28549 12764
rect 28399 12733 28411 12736
rect 28353 12727 28411 12733
rect 28537 12733 28549 12736
rect 28583 12733 28595 12767
rect 28537 12727 28595 12733
rect 28629 12767 28687 12773
rect 28629 12733 28641 12767
rect 28675 12733 28687 12767
rect 28629 12727 28687 12733
rect 27157 12699 27215 12705
rect 27157 12696 27169 12699
rect 26252 12668 27169 12696
rect 27157 12665 27169 12668
rect 27203 12665 27215 12699
rect 28644 12696 28672 12727
rect 28994 12724 29000 12776
rect 29052 12724 29058 12776
rect 30024 12773 30052 12804
rect 30834 12792 30840 12804
rect 30892 12792 30898 12844
rect 30009 12767 30067 12773
rect 30009 12733 30021 12767
rect 30055 12733 30067 12767
rect 30009 12727 30067 12733
rect 30101 12767 30159 12773
rect 30101 12733 30113 12767
rect 30147 12733 30159 12767
rect 30101 12727 30159 12733
rect 30193 12767 30251 12773
rect 30193 12733 30205 12767
rect 30239 12764 30251 12767
rect 30377 12767 30435 12773
rect 30377 12764 30389 12767
rect 30239 12736 30389 12764
rect 30239 12733 30251 12736
rect 30193 12727 30251 12733
rect 30377 12733 30389 12736
rect 30423 12733 30435 12767
rect 30377 12727 30435 12733
rect 30469 12767 30527 12773
rect 30469 12733 30481 12767
rect 30515 12764 30527 12767
rect 30653 12767 30711 12773
rect 30653 12764 30665 12767
rect 30515 12736 30665 12764
rect 30515 12733 30527 12736
rect 30469 12727 30527 12733
rect 30653 12733 30665 12736
rect 30699 12733 30711 12767
rect 30653 12727 30711 12733
rect 29089 12699 29147 12705
rect 29089 12696 29101 12699
rect 28644 12668 29101 12696
rect 27157 12659 27215 12665
rect 29089 12665 29101 12668
rect 29135 12665 29147 12699
rect 29089 12659 29147 12665
rect 29917 12699 29975 12705
rect 29917 12665 29929 12699
rect 29963 12696 29975 12699
rect 30116 12696 30144 12727
rect 29963 12668 30144 12696
rect 29963 12665 29975 12668
rect 29917 12659 29975 12665
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2832 12600 2881 12628
rect 2832 12588 2838 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 5684 12600 6101 12628
rect 5684 12588 5690 12600
rect 6089 12597 6101 12600
rect 6135 12597 6147 12631
rect 6089 12591 6147 12597
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12628 11575 12631
rect 11882 12628 11888 12640
rect 11563 12600 11888 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 15194 12588 15200 12640
rect 15252 12588 15258 12640
rect 20254 12588 20260 12640
rect 20312 12628 20318 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 20312 12600 20453 12628
rect 20312 12588 20318 12600
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 24305 12631 24363 12637
rect 24305 12597 24317 12631
rect 24351 12628 24363 12631
rect 25038 12628 25044 12640
rect 24351 12600 25044 12628
rect 24351 12597 24363 12600
rect 24305 12591 24363 12597
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 28261 12631 28319 12637
rect 28261 12597 28273 12631
rect 28307 12628 28319 12631
rect 28718 12628 28724 12640
rect 28307 12600 28724 12628
rect 28307 12597 28319 12600
rect 28261 12591 28319 12597
rect 28718 12588 28724 12600
rect 28776 12588 28782 12640
rect 552 12538 31648 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31648 12538
rect 552 12464 31648 12486
rect 4982 12384 4988 12436
rect 5040 12384 5046 12436
rect 13906 12384 13912 12436
rect 13964 12384 13970 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19484 12396 19625 12424
rect 19484 12384 19490 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 19613 12387 19671 12393
rect 21818 12384 21824 12436
rect 21876 12424 21882 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21876 12396 21925 12424
rect 21876 12384 21882 12396
rect 21913 12393 21925 12396
rect 21959 12393 21971 12427
rect 21913 12387 21971 12393
rect 26694 12384 26700 12436
rect 26752 12424 26758 12436
rect 27065 12427 27123 12433
rect 27065 12424 27077 12427
rect 26752 12396 27077 12424
rect 26752 12384 26758 12396
rect 27065 12393 27077 12396
rect 27111 12393 27123 12427
rect 27065 12387 27123 12393
rect 30834 12384 30840 12436
rect 30892 12384 30898 12436
rect 3697 12359 3755 12365
rect 3697 12356 3709 12359
rect 3528 12328 3709 12356
rect 2774 12248 2780 12300
rect 2832 12248 2838 12300
rect 3528 12297 3556 12328
rect 3697 12325 3709 12328
rect 3743 12325 3755 12359
rect 3697 12319 3755 12325
rect 9309 12359 9367 12365
rect 9309 12325 9321 12359
rect 9355 12356 9367 12359
rect 11977 12359 12035 12365
rect 11977 12356 11989 12359
rect 9355 12328 9812 12356
rect 9355 12325 9367 12328
rect 9309 12319 9367 12325
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3283 12260 3433 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 5123 12260 5273 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12288 5411 12291
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 5399 12260 5549 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3620 12220 3648 12251
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6227 12260 6377 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12288 6515 12291
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6503 12260 6653 12288
rect 6503 12257 6515 12260
rect 6457 12251 6515 12257
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6779 12260 6929 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 7055 12260 7205 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7331 12260 7481 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7607 12260 7757 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 7883 12260 8033 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8021 12257 8033 12260
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 8113 12291 8171 12297
rect 8113 12257 8125 12291
rect 8159 12288 8171 12291
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 8159 12260 8309 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12288 8447 12291
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 8435 12260 8585 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8711 12260 8861 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12288 9459 12291
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9447 12260 9597 12288
rect 9447 12257 9459 12260
rect 9401 12251 9459 12257
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 2915 12192 3648 12220
rect 8956 12220 8984 12251
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 9784 12297 9812 12328
rect 11808 12328 11989 12356
rect 11808 12297 11836 12328
rect 11977 12325 11989 12328
rect 12023 12325 12035 12359
rect 11977 12319 12035 12325
rect 14921 12359 14979 12365
rect 14921 12325 14933 12359
rect 14967 12356 14979 12359
rect 20165 12359 20223 12365
rect 14967 12328 15700 12356
rect 14967 12325 14979 12328
rect 14921 12319 14979 12325
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11563 12260 11713 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 11882 12248 11888 12300
rect 11940 12248 11946 12300
rect 13446 12248 13452 12300
rect 13504 12248 13510 12300
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13679 12260 13829 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13817 12257 13829 12260
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 15013 12291 15071 12297
rect 15013 12257 15025 12291
rect 15059 12288 15071 12291
rect 15194 12288 15200 12300
rect 15059 12260 15200 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 8956 12192 9873 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13556 12220 13584 12251
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15672 12297 15700 12328
rect 20165 12325 20177 12359
rect 20211 12356 20223 12359
rect 22189 12359 22247 12365
rect 20211 12328 20668 12356
rect 20211 12325 20223 12328
rect 20165 12319 20223 12325
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15335 12260 15485 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12257 15623 12291
rect 15565 12251 15623 12257
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 13403 12192 13584 12220
rect 15580 12220 15608 12251
rect 16298 12248 16304 12300
rect 16356 12288 16362 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16356 12260 16497 12288
rect 16356 12248 16362 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12288 16635 12291
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16623 12260 16773 12288
rect 16623 12257 16635 12260
rect 16577 12251 16635 12257
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12288 16911 12291
rect 17037 12291 17095 12297
rect 17037 12288 17049 12291
rect 16899 12260 17049 12288
rect 16899 12257 16911 12260
rect 16853 12251 16911 12257
rect 17037 12257 17049 12260
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 17175 12260 17325 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17451 12260 17601 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17727 12260 17877 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 17957 12291 18015 12297
rect 17957 12257 17969 12291
rect 18003 12288 18015 12291
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 18003 12260 18153 12288
rect 18003 12257 18015 12260
rect 17957 12251 18015 12257
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18417 12291 18475 12297
rect 18417 12288 18429 12291
rect 18279 12260 18429 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18417 12257 18429 12260
rect 18463 12257 18475 12291
rect 18417 12251 18475 12257
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 18555 12260 18705 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 18693 12257 18705 12260
rect 18739 12257 18751 12291
rect 18693 12251 18751 12257
rect 18785 12291 18843 12297
rect 18785 12257 18797 12291
rect 18831 12288 18843 12291
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18831 12260 18981 12288
rect 18831 12257 18843 12260
rect 18785 12251 18843 12257
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 19061 12291 19119 12297
rect 19061 12257 19073 12291
rect 19107 12288 19119 12291
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19107 12260 19257 12288
rect 19107 12257 19119 12260
rect 19061 12251 19119 12257
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12288 19395 12291
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 19383 12260 19533 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19521 12257 19533 12260
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 20254 12248 20260 12300
rect 20312 12248 20318 12300
rect 20640 12297 20668 12328
rect 22189 12325 22201 12359
rect 22235 12356 22247 12359
rect 30561 12359 30619 12365
rect 30561 12356 30573 12359
rect 22235 12328 22416 12356
rect 22235 12325 22247 12328
rect 22189 12319 22247 12325
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12257 20683 12291
rect 20625 12251 20683 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15580 12192 15761 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 20548 12220 20576 12251
rect 20717 12223 20775 12229
rect 20717 12220 20729 12223
rect 20548 12192 20729 12220
rect 15749 12183 15807 12189
rect 20717 12189 20729 12192
rect 20763 12189 20775 12223
rect 22020 12220 22048 12251
rect 22278 12248 22284 12300
rect 22336 12248 22342 12300
rect 22388 12297 22416 12328
rect 30116 12328 30573 12356
rect 22373 12291 22431 12297
rect 22373 12257 22385 12291
rect 22419 12257 22431 12291
rect 22373 12251 22431 12257
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 22649 12291 22707 12297
rect 22649 12288 22661 12291
rect 22511 12260 22661 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 22649 12257 22661 12260
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 24397 12291 24455 12297
rect 24397 12257 24409 12291
rect 24443 12288 24455 12291
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 24443 12260 24593 12288
rect 24443 12257 24455 12260
rect 24397 12251 24455 12257
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 24673 12291 24731 12297
rect 24673 12257 24685 12291
rect 24719 12288 24731 12291
rect 24857 12291 24915 12297
rect 24857 12288 24869 12291
rect 24719 12260 24869 12288
rect 24719 12257 24731 12260
rect 24673 12251 24731 12257
rect 24857 12257 24869 12260
rect 24903 12257 24915 12291
rect 24857 12251 24915 12257
rect 24949 12291 25007 12297
rect 24949 12257 24961 12291
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 22741 12223 22799 12229
rect 22741 12220 22753 12223
rect 22020 12192 22753 12220
rect 20717 12183 20775 12189
rect 22741 12189 22753 12192
rect 22787 12189 22799 12223
rect 24964 12220 24992 12251
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 26602 12248 26608 12300
rect 26660 12248 26666 12300
rect 26697 12291 26755 12297
rect 26697 12257 26709 12291
rect 26743 12257 26755 12291
rect 26697 12251 26755 12257
rect 26789 12291 26847 12297
rect 26789 12257 26801 12291
rect 26835 12288 26847 12291
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 26835 12260 26985 12288
rect 26835 12257 26847 12260
rect 26789 12251 26847 12257
rect 26973 12257 26985 12260
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 28353 12291 28411 12297
rect 28353 12257 28365 12291
rect 28399 12288 28411 12291
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 28399 12260 28549 12288
rect 28399 12257 28411 12260
rect 28353 12251 28411 12257
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28537 12251 28595 12257
rect 28629 12291 28687 12297
rect 28629 12257 28641 12291
rect 28675 12257 28687 12291
rect 28629 12251 28687 12257
rect 25133 12223 25191 12229
rect 25133 12220 25145 12223
rect 24964 12192 25145 12220
rect 22741 12183 22799 12189
rect 25133 12189 25145 12192
rect 25179 12189 25191 12223
rect 25133 12183 25191 12189
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12220 26571 12223
rect 26712 12220 26740 12251
rect 26559 12192 26740 12220
rect 28644 12220 28672 12251
rect 28718 12248 28724 12300
rect 28776 12248 28782 12300
rect 30116 12297 30144 12328
rect 30561 12325 30573 12328
rect 30607 12325 30619 12359
rect 30561 12319 30619 12325
rect 30101 12291 30159 12297
rect 30101 12257 30113 12291
rect 30147 12257 30159 12291
rect 30101 12251 30159 12257
rect 30374 12248 30380 12300
rect 30432 12248 30438 12300
rect 30469 12291 30527 12297
rect 30469 12257 30481 12291
rect 30515 12257 30527 12291
rect 30469 12251 30527 12257
rect 30745 12291 30803 12297
rect 30745 12257 30757 12291
rect 30791 12257 30803 12291
rect 30745 12251 30803 12257
rect 28813 12223 28871 12229
rect 28813 12220 28825 12223
rect 28644 12192 28825 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 28813 12189 28825 12192
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 30285 12223 30343 12229
rect 30285 12189 30297 12223
rect 30331 12220 30343 12223
rect 30484 12220 30512 12251
rect 30331 12192 30512 12220
rect 30331 12189 30343 12192
rect 30285 12183 30343 12189
rect 30009 12155 30067 12161
rect 30009 12121 30021 12155
rect 30055 12152 30067 12155
rect 30760 12152 30788 12251
rect 30055 12124 30788 12152
rect 30055 12121 30067 12124
rect 30009 12115 30067 12121
rect 3145 12087 3203 12093
rect 3145 12053 3157 12087
rect 3191 12084 3203 12087
rect 3234 12084 3240 12096
rect 3191 12056 3240 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 6178 12084 6184 12096
rect 6135 12056 6184 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11425 12087 11483 12093
rect 11425 12084 11437 12087
rect 11388 12056 11437 12084
rect 11388 12044 11394 12056
rect 11425 12053 11437 12056
rect 11471 12053 11483 12087
rect 11425 12047 11483 12053
rect 15102 12044 15108 12096
rect 15160 12084 15166 12096
rect 15197 12087 15255 12093
rect 15197 12084 15209 12087
rect 15160 12056 15209 12084
rect 15160 12044 15166 12056
rect 15197 12053 15209 12056
rect 15243 12053 15255 12087
rect 15197 12047 15255 12053
rect 20438 12044 20444 12096
rect 20496 12044 20502 12096
rect 24305 12087 24363 12093
rect 24305 12053 24317 12087
rect 24351 12084 24363 12087
rect 24946 12084 24952 12096
rect 24351 12056 24952 12084
rect 24351 12053 24363 12056
rect 24305 12047 24363 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 28258 12044 28264 12096
rect 28316 12044 28322 12096
rect 552 11994 31648 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31648 11994
rect 552 11920 31648 11942
rect 6270 11840 6276 11892
rect 6328 11840 6334 11892
rect 9674 11840 9680 11892
rect 9732 11840 9738 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13504 11852 13645 11880
rect 13504 11840 13510 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 16298 11840 16304 11892
rect 16356 11840 16362 11892
rect 22278 11840 22284 11892
rect 22336 11840 22342 11892
rect 26602 11840 26608 11892
rect 26660 11880 26666 11892
rect 27065 11883 27123 11889
rect 27065 11880 27077 11883
rect 26660 11852 27077 11880
rect 26660 11840 26666 11852
rect 27065 11849 27077 11852
rect 27111 11849 27123 11883
rect 27065 11843 27123 11849
rect 30374 11840 30380 11892
rect 30432 11840 30438 11892
rect 11330 11772 11336 11824
rect 11388 11772 11394 11824
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10336 11716 10517 11744
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3375 11648 3525 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3651 11648 3801 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 4065 11679 4123 11685
rect 4065 11676 4077 11679
rect 3927 11648 4077 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 4065 11645 4077 11648
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 6178 11636 6184 11688
rect 6236 11636 6242 11688
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9674 11676 9680 11688
rect 9539 11648 9680 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 10336 11685 10364 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 11348 11744 11376 11772
rect 12989 11747 13047 11753
rect 11348 11716 11468 11744
rect 10505 11707 10563 11713
rect 11440 11685 11468 11716
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13035 11716 13216 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 9769 11679 9827 11685
rect 9769 11645 9781 11679
rect 9815 11676 9827 11679
rect 9953 11679 10011 11685
rect 9953 11676 9965 11679
rect 9815 11648 9965 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 9953 11645 9965 11648
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11676 10103 11679
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 10091 11648 10241 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11645 11391 11679
rect 11333 11639 11391 11645
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11676 11575 11679
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11563 11648 11713 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11839 11648 11989 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11676 12127 11679
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 12115 11648 12265 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 9401 11611 9459 11617
rect 9401 11577 9413 11611
rect 9447 11608 9459 11611
rect 10428 11608 10456 11639
rect 9447 11580 10456 11608
rect 11348 11608 11376 11639
rect 13078 11636 13084 11688
rect 13136 11636 13142 11688
rect 13188 11685 13216 11716
rect 14016 11716 14197 11744
rect 14016 11685 14044 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 14185 11707 14243 11713
rect 20364 11716 21097 11744
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13771 11648 13921 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 12345 11611 12403 11617
rect 12345 11608 12357 11611
rect 11348 11580 12357 11608
rect 9447 11577 9459 11580
rect 9401 11571 9459 11577
rect 12345 11577 12357 11580
rect 12391 11577 12403 11611
rect 12345 11571 12403 11577
rect 13265 11611 13323 11617
rect 13265 11577 13277 11611
rect 13311 11608 13323 11611
rect 14108 11608 14136 11639
rect 15102 11636 15108 11688
rect 15160 11636 15166 11688
rect 20364 11685 20392 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 25041 11747 25099 11753
rect 25041 11744 25053 11747
rect 21085 11707 21143 11713
rect 24872 11716 25053 11744
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15243 11648 15393 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11676 15531 11679
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15519 11648 15669 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 15795 11648 15945 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 15933 11645 15945 11648
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11676 16083 11679
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 16071 11648 16221 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11645 20407 11679
rect 20349 11639 20407 11645
rect 20438 11636 20444 11688
rect 20496 11636 20502 11688
rect 24872 11685 24900 11716
rect 25041 11713 25053 11716
rect 25087 11713 25099 11747
rect 25961 11747 26019 11753
rect 25961 11744 25973 11747
rect 25041 11707 25099 11713
rect 25792 11716 25973 11744
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11676 20591 11679
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20579 11648 20729 11676
rect 20579 11645 20591 11648
rect 20533 11639 20591 11645
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20855 11648 21005 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 22557 11679 22615 11685
rect 22557 11676 22569 11679
rect 22419 11648 22569 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22557 11645 22569 11648
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 22695 11648 22845 11676
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 22925 11679 22983 11685
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 23109 11679 23167 11685
rect 23109 11676 23121 11679
rect 22971 11648 23121 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23109 11645 23121 11648
rect 23155 11645 23167 11679
rect 23109 11639 23167 11645
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11676 23259 11679
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 23247 11648 23397 11676
rect 23247 11645 23259 11648
rect 23201 11639 23259 11645
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 23937 11679 23995 11685
rect 23937 11676 23949 11679
rect 23523 11648 23949 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 23937 11645 23949 11648
rect 23983 11645 23995 11679
rect 23937 11639 23995 11645
rect 24029 11679 24087 11685
rect 24029 11645 24041 11679
rect 24075 11676 24087 11679
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 24075 11648 24225 11676
rect 24075 11645 24087 11648
rect 24029 11639 24087 11645
rect 24213 11645 24225 11648
rect 24259 11645 24271 11679
rect 24213 11639 24271 11645
rect 24305 11679 24363 11685
rect 24305 11645 24317 11679
rect 24351 11676 24363 11679
rect 24489 11679 24547 11685
rect 24489 11676 24501 11679
rect 24351 11648 24501 11676
rect 24351 11645 24363 11648
rect 24305 11639 24363 11645
rect 24489 11645 24501 11648
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 24581 11679 24639 11685
rect 24581 11645 24593 11679
rect 24627 11676 24639 11679
rect 24765 11679 24823 11685
rect 24765 11676 24777 11679
rect 24627 11648 24777 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 24765 11645 24777 11648
rect 24811 11645 24823 11679
rect 24765 11639 24823 11645
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11645 24915 11679
rect 24857 11639 24915 11645
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25792 11685 25820 11716
rect 25961 11713 25973 11716
rect 26007 11713 26019 11747
rect 25961 11707 26019 11713
rect 28169 11747 28227 11753
rect 28169 11713 28181 11747
rect 28215 11744 28227 11747
rect 30101 11747 30159 11753
rect 28215 11716 28396 11744
rect 28215 11713 28227 11716
rect 28169 11707 28227 11713
rect 25777 11679 25835 11685
rect 25777 11645 25789 11679
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 25866 11636 25872 11688
rect 25924 11636 25930 11688
rect 26145 11679 26203 11685
rect 26145 11645 26157 11679
rect 26191 11645 26203 11679
rect 26145 11639 26203 11645
rect 26237 11679 26295 11685
rect 26237 11645 26249 11679
rect 26283 11676 26295 11679
rect 26421 11679 26479 11685
rect 26421 11676 26433 11679
rect 26283 11648 26433 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 26421 11645 26433 11648
rect 26467 11645 26479 11679
rect 26421 11639 26479 11645
rect 26513 11679 26571 11685
rect 26513 11645 26525 11679
rect 26559 11676 26571 11679
rect 26697 11679 26755 11685
rect 26697 11676 26709 11679
rect 26559 11648 26709 11676
rect 26559 11645 26571 11648
rect 26513 11639 26571 11645
rect 26697 11645 26709 11648
rect 26743 11645 26755 11679
rect 26697 11639 26755 11645
rect 26789 11679 26847 11685
rect 26789 11645 26801 11679
rect 26835 11676 26847 11679
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26835 11648 26985 11676
rect 26835 11645 26847 11648
rect 26789 11639 26847 11645
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 27985 11679 28043 11685
rect 27985 11645 27997 11679
rect 28031 11645 28043 11679
rect 27985 11639 28043 11645
rect 13311 11580 14136 11608
rect 25685 11611 25743 11617
rect 13311 11577 13323 11580
rect 13265 11571 13323 11577
rect 25685 11577 25697 11611
rect 25731 11608 25743 11611
rect 26160 11608 26188 11639
rect 25731 11580 26188 11608
rect 28000 11608 28028 11639
rect 28258 11636 28264 11688
rect 28316 11636 28322 11688
rect 28368 11685 28396 11716
rect 30101 11713 30113 11747
rect 30147 11744 30159 11747
rect 30147 11716 31156 11744
rect 30147 11713 30159 11716
rect 30101 11707 30159 11713
rect 28353 11679 28411 11685
rect 28353 11645 28365 11679
rect 28399 11645 28411 11679
rect 28353 11639 28411 11645
rect 28445 11679 28503 11685
rect 28445 11645 28457 11679
rect 28491 11676 28503 11679
rect 28629 11679 28687 11685
rect 28629 11676 28641 11679
rect 28491 11648 28641 11676
rect 28491 11645 28503 11648
rect 28445 11639 28503 11645
rect 28629 11645 28641 11648
rect 28675 11645 28687 11679
rect 28629 11639 28687 11645
rect 30190 11636 30196 11688
rect 30248 11636 30254 11688
rect 31128 11685 31156 11716
rect 30469 11679 30527 11685
rect 30469 11645 30481 11679
rect 30515 11676 30527 11679
rect 30653 11679 30711 11685
rect 30653 11676 30665 11679
rect 30515 11648 30665 11676
rect 30515 11645 30527 11648
rect 30469 11639 30527 11645
rect 30653 11645 30665 11648
rect 30699 11645 30711 11679
rect 30653 11639 30711 11645
rect 30745 11679 30803 11685
rect 30745 11645 30757 11679
rect 30791 11676 30803 11679
rect 30929 11679 30987 11685
rect 30929 11676 30941 11679
rect 30791 11648 30941 11676
rect 30791 11645 30803 11648
rect 30745 11639 30803 11645
rect 30929 11645 30941 11648
rect 30975 11645 30987 11679
rect 30929 11639 30987 11645
rect 31021 11679 31079 11685
rect 31021 11645 31033 11679
rect 31067 11645 31079 11679
rect 31021 11639 31079 11645
rect 31113 11679 31171 11685
rect 31113 11645 31125 11679
rect 31159 11645 31171 11679
rect 31113 11639 31171 11645
rect 28721 11611 28779 11617
rect 28721 11608 28733 11611
rect 28000 11580 28733 11608
rect 25731 11577 25743 11580
rect 25685 11571 25743 11577
rect 28721 11577 28733 11580
rect 28767 11577 28779 11611
rect 31036 11608 31064 11639
rect 31205 11611 31263 11617
rect 31205 11608 31217 11611
rect 31036 11580 31217 11608
rect 28721 11571 28779 11577
rect 31205 11577 31217 11580
rect 31251 11577 31263 11611
rect 31205 11571 31263 11577
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 3568 11512 4169 11540
rect 3568 11500 3574 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 11241 11543 11299 11549
rect 11241 11509 11253 11543
rect 11287 11540 11299 11543
rect 11514 11540 11520 11552
rect 11287 11512 11520 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 20257 11543 20315 11549
rect 20257 11509 20269 11543
rect 20303 11540 20315 11543
rect 20898 11540 20904 11552
rect 20303 11512 20904 11540
rect 20303 11509 20315 11512
rect 20257 11503 20315 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 27893 11543 27951 11549
rect 27893 11509 27905 11543
rect 27939 11540 27951 11543
rect 28166 11540 28172 11552
rect 27939 11512 28172 11540
rect 27939 11509 27951 11512
rect 27893 11503 27951 11509
rect 28166 11500 28172 11512
rect 28224 11500 28230 11552
rect 552 11450 31648 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31648 11450
rect 552 11376 31648 11398
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7607 11308 8340 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 5261 11271 5319 11277
rect 3467 11240 3648 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 3510 11160 3516 11212
rect 3568 11160 3574 11212
rect 3620 11209 3648 11240
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5905 11271 5963 11277
rect 5307 11240 5488 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 5460 11209 5488 11240
rect 5905 11237 5917 11271
rect 5951 11268 5963 11271
rect 7837 11271 7895 11277
rect 5951 11240 6132 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11169 3663 11203
rect 3605 11163 3663 11169
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11200 3755 11203
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3743 11172 3893 11200
rect 3743 11169 3755 11172
rect 3697 11163 3755 11169
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11169 5503 11203
rect 5445 11163 5503 11169
rect 5368 11132 5396 11163
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6104 11209 6132 11240
rect 7837 11237 7849 11271
rect 7883 11268 7895 11271
rect 7883 11240 8064 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 8036 11209 8064 11240
rect 8312 11209 8340 11308
rect 9674 11296 9680 11348
rect 9732 11296 9738 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13136 11308 13277 11336
rect 13136 11296 13142 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 25866 11336 25872 11348
rect 25547 11308 25872 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 30190 11296 30196 11348
rect 30248 11336 30254 11348
rect 30653 11339 30711 11345
rect 30653 11336 30665 11339
rect 30248 11308 30665 11336
rect 30248 11296 30254 11308
rect 30653 11305 30665 11308
rect 30699 11305 30711 11339
rect 30653 11299 30711 11305
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 10060 11240 10241 11268
rect 10060 11209 10088 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 10229 11231 10287 11237
rect 13648 11240 13829 11268
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6227 11172 6377 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 6365 11163 6423 11169
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6503 11172 6653 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11200 6791 11203
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6779 11172 6929 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7055 11172 7205 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7331 11172 7481 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9815 11172 9965 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 5626 11132 5632 11144
rect 5368 11104 5632 11132
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 7944 11132 7972 11163
rect 10134 11160 10140 11212
rect 10192 11160 10198 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 13648 11209 13676 11240
rect 13817 11237 13829 11240
rect 13863 11237 13875 11271
rect 16209 11271 16267 11277
rect 16209 11268 16221 11271
rect 13817 11231 13875 11237
rect 15488 11240 16221 11268
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11655 11172 11805 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13403 11172 13553 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13541 11163 13599 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 13722 11160 13728 11212
rect 13780 11160 13786 11212
rect 15488 11209 15516 11240
rect 16209 11237 16221 11240
rect 16255 11237 16267 11271
rect 16209 11231 16267 11237
rect 17681 11271 17739 11277
rect 17681 11237 17693 11271
rect 17727 11268 17739 11271
rect 20717 11271 20775 11277
rect 20717 11268 20729 11271
rect 17727 11240 17908 11268
rect 17727 11237 17739 11240
rect 17681 11231 17739 11237
rect 17880 11209 17908 11240
rect 20548 11240 20729 11268
rect 20548 11209 20576 11240
rect 20717 11237 20729 11240
rect 20763 11237 20775 11271
rect 26053 11271 26111 11277
rect 26053 11268 26065 11271
rect 20717 11231 20775 11237
rect 25884 11240 26065 11268
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14691 11172 14841 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 14967 11172 15117 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11200 15255 11203
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 15243 11172 15393 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11169 15531 11203
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 15473 11163 15531 11169
rect 15672 11172 15853 11200
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7944 11104 8401 11132
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 15672 11064 15700 11172
rect 15841 11169 15853 11172
rect 15887 11169 15899 11203
rect 15841 11163 15899 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 17773 11203 17831 11209
rect 17773 11169 17785 11203
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 18371 11172 18521 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11200 18659 11203
rect 18785 11203 18843 11209
rect 18785 11200 18797 11203
rect 18647 11172 18797 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 18785 11169 18797 11172
rect 18831 11169 18843 11203
rect 18785 11163 18843 11169
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18923 11172 19073 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19061 11169 19073 11172
rect 19107 11169 19119 11203
rect 19061 11163 19119 11169
rect 19153 11203 19211 11209
rect 19153 11169 19165 11203
rect 19199 11200 19211 11203
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 19199 11172 19349 11200
rect 19199 11169 19211 11172
rect 19153 11163 19211 11169
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19429 11203 19487 11209
rect 19429 11169 19441 11203
rect 19475 11200 19487 11203
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19475 11172 19625 11200
rect 19475 11169 19487 11172
rect 19429 11163 19487 11169
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 19751 11172 19901 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 20027 11172 20177 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 20441 11203 20499 11209
rect 20441 11200 20453 11203
rect 20303 11172 20453 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 20441 11169 20453 11172
rect 20487 11169 20499 11203
rect 20441 11163 20499 11169
rect 20533 11203 20591 11209
rect 20533 11169 20545 11203
rect 20579 11169 20591 11203
rect 20533 11163 20591 11169
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11132 15807 11135
rect 16132 11132 16160 11163
rect 15795 11104 16160 11132
rect 17788 11132 17816 11163
rect 20622 11160 20628 11212
rect 20680 11160 20686 11212
rect 20898 11160 20904 11212
rect 20956 11160 20962 11212
rect 22830 11160 22836 11212
rect 22888 11200 22894 11212
rect 22925 11203 22983 11209
rect 22925 11200 22937 11203
rect 22888 11172 22937 11200
rect 22888 11160 22894 11172
rect 22925 11169 22937 11172
rect 22971 11169 22983 11203
rect 22925 11163 22983 11169
rect 25130 11160 25136 11212
rect 25188 11160 25194 11212
rect 25884 11209 25912 11240
rect 26053 11237 26065 11240
rect 26099 11237 26111 11271
rect 28261 11271 28319 11277
rect 28261 11268 28273 11271
rect 26053 11231 26111 11237
rect 28092 11240 28273 11268
rect 25593 11203 25651 11209
rect 25593 11169 25605 11203
rect 25639 11200 25651 11203
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 25639 11172 25789 11200
rect 25639 11169 25651 11172
rect 25593 11163 25651 11169
rect 25777 11169 25789 11172
rect 25823 11169 25835 11203
rect 25777 11163 25835 11169
rect 25869 11203 25927 11209
rect 25869 11169 25881 11203
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 25958 11160 25964 11212
rect 26016 11160 26022 11212
rect 28092 11209 28120 11240
rect 28261 11237 28273 11240
rect 28307 11237 28319 11271
rect 28261 11231 28319 11237
rect 29273 11271 29331 11277
rect 29273 11237 29285 11271
rect 29319 11268 29331 11271
rect 29319 11240 29500 11268
rect 29319 11237 29331 11240
rect 29273 11231 29331 11237
rect 27525 11203 27583 11209
rect 27525 11169 27537 11203
rect 27571 11200 27583 11203
rect 27709 11203 27767 11209
rect 27709 11200 27721 11203
rect 27571 11172 27721 11200
rect 27571 11169 27583 11172
rect 27525 11163 27583 11169
rect 27709 11169 27721 11172
rect 27755 11169 27767 11203
rect 27709 11163 27767 11169
rect 27801 11203 27859 11209
rect 27801 11169 27813 11203
rect 27847 11200 27859 11203
rect 27985 11203 28043 11209
rect 27985 11200 27997 11203
rect 27847 11172 27997 11200
rect 27847 11169 27859 11172
rect 27801 11163 27859 11169
rect 27985 11169 27997 11172
rect 28031 11169 28043 11203
rect 27985 11163 28043 11169
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11169 28135 11203
rect 28077 11163 28135 11169
rect 28166 11160 28172 11212
rect 28224 11160 28230 11212
rect 29362 11160 29368 11212
rect 29420 11160 29426 11212
rect 29472 11209 29500 11240
rect 29457 11203 29515 11209
rect 29457 11169 29469 11203
rect 29503 11169 29515 11203
rect 29457 11163 29515 11169
rect 29549 11203 29607 11209
rect 29549 11169 29561 11203
rect 29595 11200 29607 11203
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 29595 11172 29745 11200
rect 29595 11169 29607 11172
rect 29549 11163 29607 11169
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 29825 11203 29883 11209
rect 29825 11169 29837 11203
rect 29871 11200 29883 11203
rect 30009 11203 30067 11209
rect 30009 11200 30021 11203
rect 29871 11172 30021 11200
rect 29871 11169 29883 11172
rect 29825 11163 29883 11169
rect 30009 11169 30021 11172
rect 30055 11169 30067 11203
rect 30009 11163 30067 11169
rect 30101 11203 30159 11209
rect 30101 11169 30113 11203
rect 30147 11200 30159 11203
rect 30285 11203 30343 11209
rect 30285 11200 30297 11203
rect 30147 11172 30297 11200
rect 30147 11169 30159 11172
rect 30101 11163 30159 11169
rect 30285 11169 30297 11172
rect 30331 11169 30343 11203
rect 30285 11163 30343 11169
rect 30377 11203 30435 11209
rect 30377 11169 30389 11203
rect 30423 11200 30435 11203
rect 30561 11203 30619 11209
rect 30561 11200 30573 11203
rect 30423 11172 30573 11200
rect 30423 11169 30435 11172
rect 30377 11163 30435 11169
rect 30561 11169 30573 11172
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17788 11104 18245 11132
rect 15795 11101 15807 11104
rect 15749 11095 15807 11101
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 16574 11064 16580 11076
rect 15672 11036 16580 11064
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 23017 11067 23075 11073
rect 23017 11033 23029 11067
rect 23063 11064 23075 11067
rect 23842 11064 23848 11076
rect 23063 11036 23848 11064
rect 23063 11033 23075 11036
rect 23017 11027 23075 11033
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 3973 10999 4031 11005
rect 3973 10965 3985 10999
rect 4019 10996 4031 10999
rect 4062 10996 4068 11008
rect 4019 10968 4068 10996
rect 4019 10965 4031 10968
rect 3973 10959 4031 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 5537 10999 5595 11005
rect 5537 10965 5549 10999
rect 5583 10996 5595 10999
rect 5902 10996 5908 11008
rect 5583 10968 5908 10996
rect 5583 10965 5595 10968
rect 5537 10959 5595 10965
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8113 10999 8171 11005
rect 8113 10996 8125 10999
rect 8076 10968 8125 10996
rect 8076 10956 8082 10968
rect 8113 10965 8125 10968
rect 8159 10965 8171 10999
rect 8113 10959 8171 10965
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 11885 10999 11943 11005
rect 11885 10996 11897 10999
rect 11848 10968 11897 10996
rect 11848 10956 11854 10968
rect 11885 10965 11897 10968
rect 11931 10965 11943 10999
rect 11885 10959 11943 10965
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 14642 10996 14648 11008
rect 14599 10968 14648 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 17954 10956 17960 11008
rect 18012 10956 18018 11008
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 20993 10999 21051 11005
rect 20993 10996 21005 10999
rect 20772 10968 21005 10996
rect 20772 10956 20778 10968
rect 20993 10965 21005 10968
rect 21039 10965 21051 10999
rect 20993 10959 21051 10965
rect 25225 10999 25283 11005
rect 25225 10965 25237 10999
rect 25271 10996 25283 10999
rect 26050 10996 26056 11008
rect 25271 10968 26056 10996
rect 25271 10965 25283 10968
rect 25225 10959 25283 10965
rect 26050 10956 26056 10968
rect 26108 10956 26114 11008
rect 27338 10956 27344 11008
rect 27396 10996 27402 11008
rect 27433 10999 27491 11005
rect 27433 10996 27445 10999
rect 27396 10968 27445 10996
rect 27396 10956 27402 10968
rect 27433 10965 27445 10968
rect 27479 10965 27491 10999
rect 27433 10959 27491 10965
rect 552 10906 31648 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31648 10906
rect 552 10832 31648 10854
rect 5626 10752 5632 10804
rect 5684 10752 5690 10804
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6089 10795 6147 10801
rect 6089 10792 6101 10795
rect 6052 10764 6101 10792
rect 6052 10752 6058 10764
rect 6089 10761 6101 10764
rect 6135 10761 6147 10795
rect 6089 10755 6147 10761
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 10134 10792 10140 10804
rect 9539 10764 10140 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 13722 10792 13728 10804
rect 13035 10764 13728 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 16574 10752 16580 10804
rect 16632 10752 16638 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20622 10792 20628 10804
rect 20119 10764 20628 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 25869 10795 25927 10801
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 25958 10792 25964 10804
rect 25915 10764 25964 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 29362 10752 29368 10804
rect 29420 10752 29426 10804
rect 4249 10727 4307 10733
rect 4249 10724 4261 10727
rect 3528 10696 4261 10724
rect 3528 10597 3556 10696
rect 4249 10693 4261 10696
rect 4295 10693 4307 10727
rect 4249 10687 4307 10693
rect 28721 10727 28779 10733
rect 28721 10693 28733 10727
rect 28767 10724 28779 10727
rect 28767 10696 29592 10724
rect 28767 10693 28779 10696
rect 28721 10687 28779 10693
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 5077 10659 5135 10665
rect 3743 10628 3924 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 3896 10597 3924 10628
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 5123 10628 5304 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3099 10560 3433 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10557 3571 10591
rect 3513 10551 3571 10557
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10557 3939 10591
rect 3881 10551 3939 10557
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 4019 10560 4169 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4157 10557 4169 10560
rect 4203 10557 4215 10591
rect 4157 10551 4215 10557
rect 3804 10520 3832 10551
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 5276 10597 5304 10628
rect 7760 10628 8493 10656
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5399 10560 5549 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 7760 10597 7788 10628
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 16025 10659 16083 10665
rect 11747 10628 11928 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 5960 10560 6009 10588
rect 5960 10548 5966 10560
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8018 10548 8024 10600
rect 8076 10548 8082 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 4062 10520 4068 10532
rect 3804 10492 4068 10520
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 7929 10523 7987 10529
rect 7929 10489 7941 10523
rect 7975 10520 7987 10523
rect 8404 10520 8432 10551
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9907 10560 10057 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 10183 10560 10333 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10459 10560 10609 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10735 10560 10885 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 11011 10560 11161 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11425 10591 11483 10597
rect 11425 10588 11437 10591
rect 11287 10560 11437 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11425 10557 11437 10560
rect 11471 10557 11483 10591
rect 11425 10551 11483 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 7975 10492 8432 10520
rect 11532 10520 11560 10551
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 11900 10597 11928 10628
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 17589 10659 17647 10665
rect 16071 10628 16528 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10588 12035 10591
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 12023 10560 12173 10588
rect 12023 10557 12035 10560
rect 11977 10551 12035 10557
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 12161 10551 12219 10557
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10588 13139 10591
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 13127 10560 13277 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13403 10560 13829 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13955 10560 14197 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14323 10560 14565 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14642 10548 14648 10600
rect 14700 10548 14706 10600
rect 16500 10597 16528 10628
rect 17589 10625 17601 10659
rect 17635 10656 17647 10659
rect 20993 10659 21051 10665
rect 17635 10628 17816 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 16163 10560 16313 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11532 10492 12265 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 12253 10489 12265 10492
rect 12299 10489 12311 10523
rect 16408 10520 16436 10551
rect 16758 10548 16764 10600
rect 16816 10548 16822 10600
rect 17788 10597 17816 10628
rect 20993 10625 21005 10659
rect 21039 10656 21051 10659
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 21039 10628 21220 10656
rect 21039 10625 21051 10628
rect 20993 10619 21051 10625
rect 17681 10591 17739 10597
rect 17681 10557 17693 10591
rect 17727 10557 17739 10591
rect 17681 10551 17739 10557
rect 17773 10591 17831 10597
rect 17773 10557 17785 10591
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17911 10560 18061 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 20714 10588 20720 10600
rect 20211 10560 20720 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 16853 10523 16911 10529
rect 16853 10520 16865 10523
rect 16408 10492 16865 10520
rect 12253 10483 12311 10489
rect 16853 10489 16865 10492
rect 16899 10489 16911 10523
rect 17696 10520 17724 10551
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 21082 10548 21088 10600
rect 21140 10548 21146 10600
rect 21192 10597 21220 10628
rect 25976 10628 26157 10656
rect 21177 10591 21235 10597
rect 21177 10557 21189 10591
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 21315 10560 21465 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10588 21603 10591
rect 21729 10591 21787 10597
rect 21729 10588 21741 10591
rect 21591 10560 21741 10588
rect 21591 10557 21603 10560
rect 21545 10551 21603 10557
rect 21729 10557 21741 10560
rect 21775 10557 21787 10591
rect 21729 10551 21787 10557
rect 21821 10591 21879 10597
rect 21821 10557 21833 10591
rect 21867 10588 21879 10591
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 21867 10560 22017 10588
rect 21867 10557 21879 10560
rect 21821 10551 21879 10557
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10588 22155 10591
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22143 10560 22293 10588
rect 22143 10557 22155 10560
rect 22097 10551 22155 10557
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10588 22431 10591
rect 22557 10591 22615 10597
rect 22557 10588 22569 10591
rect 22419 10560 22569 10588
rect 22419 10557 22431 10560
rect 22373 10551 22431 10557
rect 22557 10557 22569 10560
rect 22603 10557 22615 10591
rect 22557 10551 22615 10557
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10588 22707 10591
rect 22833 10591 22891 10597
rect 22833 10588 22845 10591
rect 22695 10560 22845 10588
rect 22695 10557 22707 10560
rect 22649 10551 22707 10557
rect 22833 10557 22845 10560
rect 22879 10557 22891 10591
rect 22833 10551 22891 10557
rect 22925 10591 22983 10597
rect 22925 10557 22937 10591
rect 22971 10588 22983 10591
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22971 10560 23121 10588
rect 22971 10557 22983 10560
rect 22925 10551 22983 10557
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 23201 10591 23259 10597
rect 23201 10557 23213 10591
rect 23247 10588 23259 10591
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 23247 10560 23397 10588
rect 23247 10557 23259 10560
rect 23201 10551 23259 10557
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 23385 10551 23443 10557
rect 23842 10548 23848 10600
rect 23900 10548 23906 10600
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10588 23995 10591
rect 24121 10591 24179 10597
rect 24121 10588 24133 10591
rect 23983 10560 24133 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24121 10557 24133 10560
rect 24167 10557 24179 10591
rect 24121 10551 24179 10557
rect 24210 10548 24216 10600
rect 24268 10588 24274 10600
rect 24397 10591 24455 10597
rect 24397 10588 24409 10591
rect 24268 10560 24409 10588
rect 24268 10548 24274 10560
rect 24397 10557 24409 10560
rect 24443 10557 24455 10591
rect 24397 10551 24455 10557
rect 24489 10591 24547 10597
rect 24489 10557 24501 10591
rect 24535 10588 24547 10591
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24535 10560 24685 10588
rect 24535 10557 24547 10560
rect 24489 10551 24547 10557
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 24946 10548 24952 10600
rect 25004 10548 25010 10600
rect 25976 10597 26004 10628
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 29089 10659 29147 10665
rect 27295 10628 27476 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 25041 10591 25099 10597
rect 25041 10557 25053 10591
rect 25087 10588 25099 10591
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25087 10560 25237 10588
rect 25087 10557 25099 10560
rect 25041 10551 25099 10557
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 25317 10591 25375 10597
rect 25317 10557 25329 10591
rect 25363 10588 25375 10591
rect 25501 10591 25559 10597
rect 25501 10588 25513 10591
rect 25363 10560 25513 10588
rect 25363 10557 25375 10560
rect 25317 10551 25375 10557
rect 25501 10557 25513 10560
rect 25547 10557 25559 10591
rect 25501 10551 25559 10557
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 26050 10548 26056 10600
rect 26108 10548 26114 10600
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10588 26847 10591
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26835 10560 26985 10588
rect 26835 10557 26847 10560
rect 26789 10551 26847 10557
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 26973 10551 27031 10557
rect 27065 10591 27123 10597
rect 27065 10557 27077 10591
rect 27111 10557 27123 10591
rect 27065 10551 27123 10557
rect 17954 10520 17960 10532
rect 17696 10492 17960 10520
rect 16853 10483 16911 10489
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 27080 10520 27108 10551
rect 27338 10548 27344 10600
rect 27396 10548 27402 10600
rect 27448 10597 27476 10628
rect 29089 10625 29101 10659
rect 29135 10656 29147 10659
rect 29135 10628 29316 10656
rect 29135 10625 29147 10628
rect 29089 10619 29147 10625
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10557 27491 10591
rect 27433 10551 27491 10557
rect 28810 10548 28816 10600
rect 28868 10548 28874 10600
rect 29288 10597 29316 10628
rect 29564 10597 29592 10696
rect 29181 10591 29239 10597
rect 29181 10557 29193 10591
rect 29227 10557 29239 10591
rect 29181 10551 29239 10557
rect 29273 10591 29331 10597
rect 29273 10557 29285 10591
rect 29319 10557 29331 10591
rect 29273 10551 29331 10557
rect 29549 10591 29607 10597
rect 29549 10557 29561 10591
rect 29595 10557 29607 10591
rect 29549 10551 29607 10557
rect 27525 10523 27583 10529
rect 27525 10520 27537 10523
rect 27080 10492 27537 10520
rect 27525 10489 27537 10492
rect 27571 10489 27583 10523
rect 29196 10520 29224 10551
rect 29641 10523 29699 10529
rect 29641 10520 29653 10523
rect 29196 10492 29653 10520
rect 27525 10483 27583 10489
rect 29641 10489 29653 10492
rect 29687 10489 29699 10523
rect 29641 10483 29699 10489
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3234 10452 3240 10464
rect 3007 10424 3240 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 7650 10412 7656 10464
rect 7708 10412 7714 10464
rect 9766 10412 9772 10464
rect 9824 10412 9830 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 17920 10424 18153 10452
rect 17920 10412 17926 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 22922 10412 22928 10464
rect 22980 10452 22986 10464
rect 23477 10455 23535 10461
rect 23477 10452 23489 10455
rect 22980 10424 23489 10452
rect 22980 10412 22986 10424
rect 23477 10421 23489 10424
rect 23523 10421 23535 10455
rect 23477 10415 23535 10421
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 24213 10455 24271 10461
rect 24213 10452 24225 10455
rect 23716 10424 24225 10452
rect 23716 10412 23722 10424
rect 24213 10421 24225 10424
rect 24259 10421 24271 10455
rect 24213 10415 24271 10421
rect 24762 10412 24768 10464
rect 24820 10412 24826 10464
rect 25222 10412 25228 10464
rect 25280 10452 25286 10464
rect 25593 10455 25651 10461
rect 25593 10452 25605 10455
rect 25280 10424 25605 10452
rect 25280 10412 25286 10424
rect 25593 10421 25605 10424
rect 25639 10421 25651 10455
rect 25593 10415 25651 10421
rect 26694 10412 26700 10464
rect 26752 10412 26758 10464
rect 552 10362 31648 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31648 10362
rect 552 10288 31648 10310
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 5224 10220 5365 10248
rect 5224 10208 5230 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5353 10211 5411 10217
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 7515 10220 8524 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 3881 10183 3939 10189
rect 3881 10180 3893 10183
rect 3160 10152 3893 10180
rect 3160 10121 3188 10152
rect 3881 10149 3893 10152
rect 3927 10149 3939 10183
rect 5905 10183 5963 10189
rect 5905 10180 5917 10183
rect 3881 10143 3939 10149
rect 5460 10152 5917 10180
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 3234 10072 3240 10124
rect 3292 10072 3298 10124
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3375 10084 3525 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3651 10084 3801 10112
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 5460 10121 5488 10152
rect 5905 10149 5917 10152
rect 5951 10149 5963 10183
rect 5905 10143 5963 10149
rect 7745 10183 7803 10189
rect 7745 10149 7757 10183
rect 7791 10180 7803 10183
rect 7791 10152 8248 10180
rect 7791 10149 7803 10152
rect 7745 10143 7803 10149
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 5000 10084 5181 10112
rect 5000 9976 5028 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 7561 10115 7619 10121
rect 6135 10084 6316 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5828 10044 5856 10075
rect 5123 10016 5856 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 6181 9979 6239 9985
rect 6181 9976 6193 9979
rect 5000 9948 6193 9976
rect 6181 9945 6193 9948
rect 6227 9945 6239 9979
rect 6181 9939 6239 9945
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 3234 9908 3240 9920
rect 3099 9880 3240 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 6288 9908 6316 10084
rect 7561 10081 7573 10115
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7576 10044 7604 10075
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 8220 10121 8248 10152
rect 8496 10121 8524 10220
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9640 10220 9873 10248
rect 9640 10208 9646 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 16393 10251 16451 10257
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 16758 10248 16764 10260
rect 16439 10220 16764 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 21082 10208 21088 10260
rect 21140 10248 21146 10260
rect 21637 10251 21695 10257
rect 21637 10248 21649 10251
rect 21140 10220 21649 10248
rect 21140 10208 21146 10220
rect 21637 10217 21649 10220
rect 21683 10217 21695 10251
rect 21637 10211 21695 10217
rect 22830 10208 22836 10260
rect 22888 10208 22894 10260
rect 23569 10251 23627 10257
rect 23569 10217 23581 10251
rect 23615 10248 23627 10251
rect 24210 10248 24216 10260
rect 23615 10220 24216 10248
rect 23615 10217 23627 10220
rect 23569 10211 23627 10217
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 24397 10251 24455 10257
rect 24397 10217 24409 10251
rect 24443 10248 24455 10251
rect 24946 10248 24952 10260
rect 24443 10220 24952 10248
rect 24443 10217 24455 10220
rect 24397 10211 24455 10217
rect 24946 10208 24952 10220
rect 25004 10208 25010 10260
rect 25130 10208 25136 10260
rect 25188 10208 25194 10260
rect 28810 10208 28816 10260
rect 28868 10208 28874 10260
rect 16945 10183 17003 10189
rect 16945 10180 16957 10183
rect 16776 10152 16957 10180
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 8128 10044 8156 10075
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 16776 10121 16804 10152
rect 16945 10149 16957 10152
rect 16991 10149 17003 10183
rect 24762 10180 24768 10192
rect 16945 10143 17003 10149
rect 24228 10152 24768 10180
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10112 16543 10115
rect 16669 10115 16727 10121
rect 16669 10112 16681 10115
rect 16531 10084 16681 10112
rect 16531 10081 16543 10084
rect 16485 10075 16543 10081
rect 16669 10081 16681 10084
rect 16715 10081 16727 10115
rect 16669 10075 16727 10081
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 17862 10072 17868 10124
rect 17920 10072 17926 10124
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18095 10084 18245 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18371 10084 18521 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 8573 10047 8631 10053
rect 8573 10044 8585 10047
rect 7576 10016 7696 10044
rect 8128 10016 8585 10044
rect 7668 9976 7696 10016
rect 8573 10013 8585 10016
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 17972 10044 18000 10075
rect 19794 10072 19800 10124
rect 19852 10072 19858 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10081 19947 10115
rect 19889 10075 19947 10081
rect 19981 10115 20039 10121
rect 19981 10081 19993 10115
rect 20027 10112 20039 10115
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 20027 10084 20177 10112
rect 20027 10081 20039 10084
rect 19981 10075 20039 10081
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20165 10075 20223 10081
rect 20257 10115 20315 10121
rect 20257 10081 20269 10115
rect 20303 10112 20315 10115
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 20303 10084 20453 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 20441 10081 20453 10084
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 20717 10115 20775 10121
rect 20717 10112 20729 10115
rect 20579 10084 20729 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 20717 10081 20729 10084
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 20809 10115 20867 10121
rect 20809 10081 20821 10115
rect 20855 10112 20867 10115
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 20855 10084 21281 10112
rect 20855 10081 20867 10084
rect 20809 10075 20867 10081
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 21407 10084 21557 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 21545 10081 21557 10084
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 17819 10016 18000 10044
rect 19705 10047 19763 10053
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 19904 10044 19932 10075
rect 22922 10072 22928 10124
rect 22980 10072 22986 10124
rect 23658 10072 23664 10124
rect 23716 10072 23722 10124
rect 24228 10121 24256 10152
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 27341 10183 27399 10189
rect 27341 10180 27353 10183
rect 26620 10152 27353 10180
rect 24213 10115 24271 10121
rect 24213 10081 24225 10115
rect 24259 10081 24271 10115
rect 24213 10075 24271 10081
rect 24305 10115 24363 10121
rect 24305 10081 24317 10115
rect 24351 10081 24363 10115
rect 24305 10075 24363 10081
rect 19751 10016 19932 10044
rect 24121 10047 24179 10053
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 24121 10013 24133 10047
rect 24167 10044 24179 10047
rect 24320 10044 24348 10075
rect 25222 10072 25228 10124
rect 25280 10072 25286 10124
rect 26620 10121 26648 10152
rect 27341 10149 27353 10152
rect 27387 10149 27399 10183
rect 29641 10183 29699 10189
rect 29641 10180 29653 10183
rect 27341 10143 27399 10149
rect 29472 10152 29653 10180
rect 26605 10115 26663 10121
rect 26605 10081 26617 10115
rect 26651 10081 26663 10115
rect 26605 10075 26663 10081
rect 26694 10072 26700 10124
rect 26752 10072 26758 10124
rect 29472 10121 29500 10152
rect 29641 10149 29653 10152
rect 29687 10149 29699 10183
rect 29641 10143 29699 10149
rect 26789 10115 26847 10121
rect 26789 10081 26801 10115
rect 26835 10112 26847 10115
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26835 10084 26985 10112
rect 26835 10081 26847 10084
rect 26789 10075 26847 10081
rect 26973 10081 26985 10084
rect 27019 10081 27031 10115
rect 26973 10075 27031 10081
rect 27065 10115 27123 10121
rect 27065 10081 27077 10115
rect 27111 10112 27123 10115
rect 27249 10115 27307 10121
rect 27249 10112 27261 10115
rect 27111 10084 27261 10112
rect 27111 10081 27123 10084
rect 27065 10075 27123 10081
rect 27249 10081 27261 10084
rect 27295 10081 27307 10115
rect 27249 10075 27307 10081
rect 28905 10115 28963 10121
rect 28905 10081 28917 10115
rect 28951 10112 28963 10115
rect 29089 10115 29147 10121
rect 29089 10112 29101 10115
rect 28951 10084 29101 10112
rect 28951 10081 28963 10084
rect 28905 10075 28963 10081
rect 29089 10081 29101 10084
rect 29135 10081 29147 10115
rect 29089 10075 29147 10081
rect 29181 10115 29239 10121
rect 29181 10081 29193 10115
rect 29227 10112 29239 10115
rect 29365 10115 29423 10121
rect 29365 10112 29377 10115
rect 29227 10084 29377 10112
rect 29227 10081 29239 10084
rect 29181 10075 29239 10081
rect 29365 10081 29377 10084
rect 29411 10081 29423 10115
rect 29365 10075 29423 10081
rect 29457 10115 29515 10121
rect 29457 10081 29469 10115
rect 29503 10081 29515 10115
rect 29457 10075 29515 10081
rect 29546 10072 29552 10124
rect 29604 10072 29610 10124
rect 24167 10016 24348 10044
rect 24167 10013 24179 10016
rect 24121 10007 24179 10013
rect 8297 9979 8355 9985
rect 8297 9976 8309 9979
rect 7668 9948 8309 9976
rect 8297 9945 8309 9948
rect 8343 9945 8355 9979
rect 8297 9939 8355 9945
rect 4847 9880 6316 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8021 9911 8079 9917
rect 8021 9908 8033 9911
rect 7984 9880 8033 9908
rect 7984 9868 7990 9880
rect 8021 9877 8033 9880
rect 8067 9877 8079 9911
rect 8021 9871 8079 9877
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18601 9911 18659 9917
rect 18601 9908 18613 9911
rect 18472 9880 18613 9908
rect 18472 9868 18478 9880
rect 18601 9877 18613 9880
rect 18647 9877 18659 9911
rect 18601 9871 18659 9877
rect 26513 9911 26571 9917
rect 26513 9877 26525 9911
rect 26559 9908 26571 9911
rect 26602 9908 26608 9920
rect 26559 9880 26608 9908
rect 26559 9877 26571 9880
rect 26513 9871 26571 9877
rect 26602 9868 26608 9880
rect 26660 9868 26666 9920
rect 552 9818 31648 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31648 9818
rect 552 9744 31648 9766
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5169 9707 5227 9713
rect 5169 9704 5181 9707
rect 4948 9676 5181 9704
rect 4948 9664 4954 9676
rect 5169 9673 5181 9676
rect 5215 9673 5227 9707
rect 5169 9667 5227 9673
rect 16669 9707 16727 9713
rect 16669 9673 16681 9707
rect 16715 9704 16727 9707
rect 16850 9704 16856 9716
rect 16715 9676 16856 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 20165 9707 20223 9713
rect 20165 9704 20177 9707
rect 19852 9676 20177 9704
rect 19852 9664 19858 9676
rect 20165 9673 20177 9676
rect 20211 9673 20223 9707
rect 20165 9667 20223 9673
rect 29089 9707 29147 9713
rect 29089 9673 29101 9707
rect 29135 9704 29147 9707
rect 29546 9704 29552 9716
rect 29135 9676 29552 9704
rect 29135 9673 29147 9676
rect 29089 9667 29147 9673
rect 29546 9664 29552 9676
rect 29604 9664 29610 9716
rect 15105 9639 15163 9645
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 15151 9608 15608 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 10965 9571 11023 9577
rect 4939 9540 5396 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3375 9472 3525 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3651 9472 3801 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3927 9472 4077 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4706 9500 4712 9512
rect 4571 9472 4712 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5368 9509 5396 9540
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 14829 9571 14887 9577
rect 11011 9540 11560 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 4617 9435 4675 9441
rect 4617 9401 4629 9435
rect 4663 9432 4675 9435
rect 4816 9432 4844 9463
rect 4663 9404 4844 9432
rect 5276 9432 5304 9463
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5276 9404 5457 9432
rect 4663 9401 4675 9404
rect 4617 9395 4675 9401
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 5445 9395 5503 9401
rect 7837 9435 7895 9441
rect 7837 9401 7849 9435
rect 7883 9432 7895 9435
rect 8036 9432 8064 9463
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 11532 9509 11560 9540
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 14875 9540 15332 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8803 9472 8953 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9079 9472 9229 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 9355 9472 9505 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9631 9472 9781 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9907 9472 10057 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 10183 9472 10333 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 10597 9503 10655 9509
rect 10597 9500 10609 9503
rect 10459 9472 10609 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 10597 9469 10609 9472
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10735 9472 10885 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9469 11483 9503
rect 11425 9463 11483 9469
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 7883 9404 8064 9432
rect 8481 9435 8539 9441
rect 7883 9401 7895 9404
rect 7837 9395 7895 9401
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8680 9432 8708 9463
rect 8527 9404 8708 9432
rect 11440 9432 11468 9463
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 15304 9509 15332 9540
rect 15580 9509 15608 9608
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 28721 9571 28779 9577
rect 18371 9540 18736 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 13035 9472 13185 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13173 9469 13185 9472
rect 13219 9469 13231 9503
rect 13173 9463 13231 9469
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9500 13323 9503
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13311 9472 13645 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13771 9472 13921 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14047 9472 14197 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14323 9472 14473 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14599 9472 14749 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15565 9463 15623 9469
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9500 16819 9503
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16807 9472 16957 9500
rect 16807 9469 16819 9472
rect 16761 9463 16819 9469
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17037 9503 17095 9509
rect 17037 9469 17049 9503
rect 17083 9500 17095 9503
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 17083 9472 17233 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 11609 9435 11667 9441
rect 11609 9432 11621 9435
rect 11440 9404 11621 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 11609 9401 11621 9404
rect 11655 9401 11667 9435
rect 11609 9395 11667 9401
rect 12713 9435 12771 9441
rect 12713 9401 12725 9435
rect 12759 9432 12771 9435
rect 12912 9432 12940 9463
rect 12759 9404 12940 9432
rect 15212 9432 15240 9463
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 15212 9404 15393 9432
rect 12759 9401 12771 9404
rect 12713 9395 12771 9401
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 17328 9432 17356 9463
rect 17402 9460 17408 9512
rect 17460 9460 17466 9512
rect 18414 9460 18420 9512
rect 18472 9460 18478 9512
rect 18708 9509 18736 9540
rect 28721 9537 28733 9571
rect 28767 9568 28779 9571
rect 28767 9540 29592 9568
rect 28767 9537 28779 9540
rect 28721 9531 28779 9537
rect 18693 9503 18751 9509
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 18785 9503 18843 9509
rect 18785 9469 18797 9503
rect 18831 9500 18843 9503
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18831 9472 18981 9500
rect 18831 9469 18843 9472
rect 18785 9463 18843 9469
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9500 19119 9503
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 19107 9472 19257 9500
rect 19107 9469 19119 9472
rect 19061 9463 19119 9469
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9500 19395 9503
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19383 9472 19533 9500
rect 19383 9469 19395 9472
rect 19337 9463 19395 9469
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19659 9472 19809 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19935 9472 20085 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 22465 9503 22523 9509
rect 22465 9500 22477 9503
rect 22327 9472 22477 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 22465 9469 22477 9472
rect 22511 9469 22523 9503
rect 22465 9463 22523 9469
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9500 22615 9503
rect 22741 9503 22799 9509
rect 22741 9500 22753 9503
rect 22603 9472 22753 9500
rect 22603 9469 22615 9472
rect 22557 9463 22615 9469
rect 22741 9469 22753 9472
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 22833 9503 22891 9509
rect 22833 9469 22845 9503
rect 22879 9500 22891 9503
rect 23017 9503 23075 9509
rect 23017 9500 23029 9503
rect 22879 9472 23029 9500
rect 22879 9469 22891 9472
rect 22833 9463 22891 9469
rect 23017 9469 23029 9472
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9469 23167 9503
rect 23109 9463 23167 9469
rect 17497 9435 17555 9441
rect 17497 9432 17509 9435
rect 17328 9404 17509 9432
rect 15381 9395 15439 9401
rect 17497 9401 17509 9404
rect 17543 9401 17555 9435
rect 23124 9432 23152 9463
rect 23198 9460 23204 9512
rect 23256 9460 23262 9512
rect 26513 9503 26571 9509
rect 26513 9469 26525 9503
rect 26559 9469 26571 9503
rect 26513 9463 26571 9469
rect 23293 9435 23351 9441
rect 23293 9432 23305 9435
rect 23124 9404 23305 9432
rect 17497 9395 17555 9401
rect 23293 9401 23305 9404
rect 23339 9401 23351 9435
rect 26528 9432 26556 9463
rect 26602 9460 26608 9512
rect 26660 9460 26666 9512
rect 26697 9503 26755 9509
rect 26697 9469 26709 9503
rect 26743 9500 26755 9503
rect 26881 9503 26939 9509
rect 26881 9500 26893 9503
rect 26743 9472 26893 9500
rect 26743 9469 26755 9472
rect 26697 9463 26755 9469
rect 26881 9469 26893 9472
rect 26927 9469 26939 9503
rect 26881 9463 26939 9469
rect 26973 9503 27031 9509
rect 26973 9469 26985 9503
rect 27019 9500 27031 9503
rect 27157 9503 27215 9509
rect 27157 9500 27169 9503
rect 27019 9472 27169 9500
rect 27019 9469 27031 9472
rect 26973 9463 27031 9469
rect 27157 9469 27169 9472
rect 27203 9469 27215 9503
rect 27157 9463 27215 9469
rect 28810 9460 28816 9512
rect 28868 9460 28874 9512
rect 29564 9509 29592 9540
rect 29181 9503 29239 9509
rect 29181 9469 29193 9503
rect 29227 9500 29239 9503
rect 29365 9503 29423 9509
rect 29365 9500 29377 9503
rect 29227 9472 29377 9500
rect 29227 9469 29239 9472
rect 29181 9463 29239 9469
rect 29365 9469 29377 9472
rect 29411 9469 29423 9503
rect 29365 9463 29423 9469
rect 29457 9503 29515 9509
rect 29457 9469 29469 9503
rect 29503 9469 29515 9503
rect 29457 9463 29515 9469
rect 29549 9503 29607 9509
rect 29549 9469 29561 9503
rect 29595 9469 29607 9503
rect 29549 9463 29607 9469
rect 27249 9435 27307 9441
rect 27249 9432 27261 9435
rect 26528 9404 27261 9432
rect 23293 9395 23351 9401
rect 27249 9401 27261 9404
rect 27295 9401 27307 9435
rect 29472 9432 29500 9463
rect 29641 9435 29699 9441
rect 29641 9432 29653 9435
rect 29472 9404 29653 9432
rect 27249 9395 27307 9401
rect 29641 9401 29653 9404
rect 29687 9401 29699 9435
rect 29641 9395 29699 9401
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3660 9336 4169 9364
rect 3660 9324 3666 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4157 9327 4215 9333
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8570 9364 8576 9376
rect 8159 9336 8576 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15344 9336 15669 9364
rect 15344 9324 15350 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 15657 9327 15715 9333
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 22646 9364 22652 9376
rect 22235 9336 22652 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 26421 9367 26479 9373
rect 26421 9333 26433 9367
rect 26467 9364 26479 9367
rect 26510 9364 26516 9376
rect 26467 9336 26516 9364
rect 26467 9333 26479 9336
rect 26421 9327 26479 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 552 9274 31648 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31648 9274
rect 552 9200 31648 9222
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4706 9160 4712 9172
rect 4571 9132 4712 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 8662 9120 8668 9172
rect 8720 9120 8726 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12860 9132 13001 9160
rect 12860 9120 12866 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 17129 9163 17187 9169
rect 17129 9129 17141 9163
rect 17175 9160 17187 9163
rect 17402 9160 17408 9172
rect 17175 9132 17408 9160
rect 17175 9129 17187 9132
rect 17129 9123 17187 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 23198 9120 23204 9172
rect 23256 9120 23262 9172
rect 28810 9120 28816 9172
rect 28868 9120 28874 9172
rect 4801 9095 4859 9101
rect 4801 9092 4813 9095
rect 4356 9064 4813 9092
rect 3602 8984 3608 9036
rect 3660 8984 3666 9036
rect 4356 9033 4384 9064
rect 4801 9061 4813 9064
rect 4847 9061 4859 9095
rect 4801 9055 4859 9061
rect 12621 9095 12679 9101
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 15197 9095 15255 9101
rect 12667 9064 13216 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 3697 9027 3755 9033
rect 3697 8993 3709 9027
rect 3743 8993 3755 9027
rect 3697 8987 3755 8993
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 4433 8987 4491 8993
rect 4540 8996 4721 9024
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 3712 8956 3740 8987
rect 3559 8928 3740 8956
rect 4249 8959 4307 8965
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4448 8956 4476 8987
rect 4295 8928 4476 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 3789 8891 3847 8897
rect 3789 8857 3801 8891
rect 3835 8888 3847 8891
rect 4540 8888 4568 8996
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 7558 9024 7564 9036
rect 7515 8996 7564 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8570 8984 8576 9036
rect 8628 8984 8634 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 13188 9033 13216 9064
rect 15197 9061 15209 9095
rect 15243 9092 15255 9095
rect 29641 9095 29699 9101
rect 29641 9092 29653 9095
rect 15243 9064 15424 9092
rect 15243 9061 15255 9064
rect 15197 9055 15255 9061
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11204 8996 11345 9024
rect 11204 8984 11210 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 9024 11575 9027
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11563 8996 11713 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11839 8996 11989 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12253 9027 12311 9033
rect 12253 9024 12265 9027
rect 12115 8996 12265 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12253 8993 12265 8996
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12391 8996 12541 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 15013 9027 15071 9033
rect 15013 8993 15025 9027
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11440 8956 11468 8987
rect 11287 8928 11468 8956
rect 13096 8956 13124 8987
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 13096 8928 13277 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 15028 8956 15056 8987
rect 15286 8984 15292 9036
rect 15344 8984 15350 9036
rect 15396 9033 15424 9064
rect 29472 9064 29653 9092
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15519 8996 15669 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 17221 9027 17279 9033
rect 17221 8993 17233 9027
rect 17267 9024 17279 9027
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17267 8996 17417 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 17497 9027 17555 9033
rect 17497 8993 17509 9027
rect 17543 9024 17555 9027
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 17543 8996 17693 9024
rect 17543 8993 17555 8996
rect 17497 8987 17555 8993
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15028 8928 15761 8956
rect 13265 8919 13323 8925
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 17788 8956 17816 8987
rect 17862 8984 17868 9036
rect 17920 8984 17926 9036
rect 19058 8984 19064 9036
rect 19116 8984 19122 9036
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 9024 19579 9027
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 19567 8996 19717 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 19705 8993 19717 8996
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 9024 19855 9027
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19843 8996 19993 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 19981 8993 19993 8996
rect 20027 8993 20039 9027
rect 19981 8987 20039 8993
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 20119 8996 20269 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 20395 8996 20545 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 20533 8993 20545 8996
rect 20579 8993 20591 9027
rect 20533 8987 20591 8993
rect 20625 9027 20683 9033
rect 20625 8993 20637 9027
rect 20671 9024 20683 9027
rect 20809 9027 20867 9033
rect 20809 9024 20821 9027
rect 20671 8996 20821 9024
rect 20671 8993 20683 8996
rect 20625 8987 20683 8993
rect 20809 8993 20821 8996
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21361 9027 21419 9033
rect 21361 9024 21373 9027
rect 20947 8996 21373 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 21361 8993 21373 8996
rect 21407 8993 21419 9027
rect 21361 8987 21419 8993
rect 21453 9027 21511 9033
rect 21453 8993 21465 9027
rect 21499 9024 21511 9027
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 21499 8996 21649 9024
rect 21499 8993 21511 8996
rect 21453 8987 21511 8993
rect 21637 8993 21649 8996
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 21729 9027 21787 9033
rect 21729 8993 21741 9027
rect 21775 9024 21787 9027
rect 21913 9027 21971 9033
rect 21913 9024 21925 9027
rect 21775 8996 21925 9024
rect 21775 8993 21787 8996
rect 21729 8987 21787 8993
rect 21913 8993 21925 8996
rect 21959 8993 21971 9027
rect 21913 8987 21971 8993
rect 22005 9027 22063 9033
rect 22005 8993 22017 9027
rect 22051 9024 22063 9027
rect 22189 9027 22247 9033
rect 22189 9024 22201 9027
rect 22051 8996 22201 9024
rect 22051 8993 22063 8996
rect 22005 8987 22063 8993
rect 22189 8993 22201 8996
rect 22235 8993 22247 9027
rect 22189 8987 22247 8993
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17788 8928 17969 8956
rect 15749 8919 15807 8925
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 22296 8956 22324 8987
rect 22370 8984 22376 9036
rect 22428 8984 22434 9036
rect 22646 8984 22652 9036
rect 22704 8984 22710 9036
rect 23293 9027 23351 9033
rect 23293 8993 23305 9027
rect 23339 9024 23351 9027
rect 23477 9027 23535 9033
rect 23477 9024 23489 9027
rect 23339 8996 23489 9024
rect 23339 8993 23351 8996
rect 23293 8987 23351 8993
rect 23477 8993 23489 8996
rect 23523 8993 23535 9027
rect 23477 8987 23535 8993
rect 23569 9027 23627 9033
rect 23569 8993 23581 9027
rect 23615 9024 23627 9027
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 23615 8996 23765 9024
rect 23615 8993 23627 8996
rect 23569 8987 23627 8993
rect 23753 8993 23765 8996
rect 23799 8993 23811 9027
rect 23753 8987 23811 8993
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24029 9027 24087 9033
rect 24029 9024 24041 9027
rect 23891 8996 24041 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24029 8993 24041 8996
rect 24075 8993 24087 9027
rect 24029 8987 24087 8993
rect 24121 9027 24179 9033
rect 24121 8993 24133 9027
rect 24167 9024 24179 9027
rect 24305 9027 24363 9033
rect 24305 9024 24317 9027
rect 24167 8996 24317 9024
rect 24167 8993 24179 8996
rect 24121 8987 24179 8993
rect 24305 8993 24317 8996
rect 24351 8993 24363 9027
rect 24305 8987 24363 8993
rect 24397 9027 24455 9033
rect 24397 8993 24409 9027
rect 24443 8993 24455 9027
rect 24397 8987 24455 8993
rect 22465 8959 22523 8965
rect 22465 8956 22477 8959
rect 22296 8928 22477 8956
rect 17957 8919 18015 8925
rect 22465 8925 22477 8928
rect 22511 8925 22523 8959
rect 24412 8956 24440 8987
rect 24486 8984 24492 9036
rect 24544 8984 24550 9036
rect 26510 8984 26516 9036
rect 26568 8984 26574 9036
rect 29472 9033 29500 9064
rect 29641 9061 29653 9064
rect 29687 9061 29699 9095
rect 29641 9055 29699 9061
rect 26605 9027 26663 9033
rect 26605 8993 26617 9027
rect 26651 9024 26663 9027
rect 26789 9027 26847 9033
rect 26789 9024 26801 9027
rect 26651 8996 26801 9024
rect 26651 8993 26663 8996
rect 26605 8987 26663 8993
rect 26789 8993 26801 8996
rect 26835 8993 26847 9027
rect 26789 8987 26847 8993
rect 26881 9027 26939 9033
rect 26881 8993 26893 9027
rect 26927 9024 26939 9027
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 26927 8996 27077 9024
rect 26927 8993 26939 8996
rect 26881 8987 26939 8993
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27065 8987 27123 8993
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 9024 28963 9027
rect 29089 9027 29147 9033
rect 29089 9024 29101 9027
rect 28951 8996 29101 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 29089 8993 29101 8996
rect 29135 8993 29147 9027
rect 29089 8987 29147 8993
rect 29181 9027 29239 9033
rect 29181 8993 29193 9027
rect 29227 9024 29239 9027
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 29227 8996 29377 9024
rect 29227 8993 29239 8996
rect 29181 8987 29239 8993
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 29365 8987 29423 8993
rect 29457 9027 29515 9033
rect 29457 8993 29469 9027
rect 29503 8993 29515 9027
rect 29457 8987 29515 8993
rect 29546 8984 29552 9036
rect 29604 8984 29610 9036
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24412 8928 24593 8956
rect 22465 8919 22523 8925
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 3835 8860 4568 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 8018 8820 8024 8832
rect 7607 8792 8024 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15102 8820 15108 8832
rect 14967 8792 15108 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 18966 8780 18972 8832
rect 19024 8780 19030 8832
rect 19429 8823 19487 8829
rect 19429 8789 19441 8823
rect 19475 8820 19487 8823
rect 19610 8820 19616 8832
rect 19475 8792 19616 8820
rect 19475 8789 19487 8792
rect 19429 8783 19487 8789
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 22741 8823 22799 8829
rect 22741 8820 22753 8823
rect 21968 8792 22753 8820
rect 21968 8780 21974 8792
rect 22741 8789 22753 8792
rect 22787 8789 22799 8823
rect 22741 8783 22799 8789
rect 26694 8780 26700 8832
rect 26752 8820 26758 8832
rect 27157 8823 27215 8829
rect 27157 8820 27169 8823
rect 26752 8792 27169 8820
rect 26752 8780 26758 8792
rect 27157 8789 27169 8792
rect 27203 8789 27215 8823
rect 27157 8783 27215 8789
rect 552 8730 31648 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31648 8730
rect 552 8656 31648 8678
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11204 8588 11529 8616
rect 11204 8576 11210 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8616 17279 8619
rect 17862 8616 17868 8628
rect 17267 8588 17868 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18969 8619 19027 8625
rect 18969 8585 18981 8619
rect 19015 8616 19027 8619
rect 19058 8616 19064 8628
rect 19015 8588 19064 8616
rect 19015 8585 19027 8588
rect 18969 8579 19027 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 22370 8616 22376 8628
rect 21867 8588 22376 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 24029 8619 24087 8625
rect 24029 8585 24041 8619
rect 24075 8616 24087 8619
rect 24486 8616 24492 8628
rect 24075 8588 24492 8616
rect 24075 8585 24087 8588
rect 24029 8579 24087 8585
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 29365 8619 29423 8625
rect 29365 8585 29377 8619
rect 29411 8616 29423 8619
rect 29546 8616 29552 8628
rect 29411 8588 29552 8616
rect 29411 8585 29423 8588
rect 29365 8579 29423 8585
rect 29546 8576 29552 8588
rect 29604 8576 29610 8628
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 19076 8520 19809 8548
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 16991 8452 17724 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 7374 8372 7380 8424
rect 7432 8372 7438 8424
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 7699 8384 7849 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 7837 8375 7895 8381
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 7975 8384 8125 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 8113 8381 8125 8384
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8478 8412 8484 8424
rect 8251 8384 8484 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8662 8372 8668 8424
rect 8720 8372 8726 8424
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8987 8384 9137 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9263 8384 9413 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9539 8384 9689 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9677 8381 9689 8384
rect 9723 8381 9735 8415
rect 9677 8375 9735 8381
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9815 8384 9965 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9953 8381 9965 8384
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 10091 8384 10241 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 10229 8381 10241 8384
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 10367 8384 10517 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 10612 8344 10640 8375
rect 10686 8372 10692 8424
rect 10744 8372 10750 8424
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 11388 8384 11437 8412
rect 11388 8372 11394 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 15102 8372 15108 8424
rect 15160 8372 15166 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15243 8384 15393 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15519 8384 15669 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15795 8384 15945 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 17034 8372 17040 8424
rect 17092 8372 17098 8424
rect 17696 8421 17724 8452
rect 19076 8421 19104 8520
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 19610 8480 19616 8492
rect 19352 8452 19616 8480
rect 19352 8421 19380 8452
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 17359 8384 17509 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17589 8415 17647 8421
rect 17589 8381 17601 8415
rect 17635 8381 17647 8415
rect 17589 8375 17647 8381
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8381 17739 8415
rect 17681 8375 17739 8381
rect 19061 8415 19119 8421
rect 19061 8381 19073 8415
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8412 19579 8415
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19567 8384 19717 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 10781 8347 10839 8353
rect 10781 8344 10793 8347
rect 10612 8316 10793 8344
rect 10781 8313 10793 8316
rect 10827 8313 10839 8347
rect 17604 8344 17632 8375
rect 17773 8347 17831 8353
rect 17773 8344 17785 8347
rect 17604 8316 17785 8344
rect 10781 8307 10839 8313
rect 17773 8313 17785 8316
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8344 19303 8347
rect 19444 8344 19472 8375
rect 21910 8372 21916 8424
rect 21968 8372 21974 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8412 24179 8415
rect 24305 8415 24363 8421
rect 24305 8412 24317 8415
rect 24167 8384 24317 8412
rect 24167 8381 24179 8384
rect 24121 8375 24179 8381
rect 24305 8381 24317 8384
rect 24351 8381 24363 8415
rect 24305 8375 24363 8381
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 19291 8316 19472 8344
rect 24412 8344 24440 8375
rect 24486 8372 24492 8424
rect 24544 8372 24550 8424
rect 26694 8372 26700 8424
rect 26752 8372 26758 8424
rect 26789 8415 26847 8421
rect 26789 8381 26801 8415
rect 26835 8381 26847 8415
rect 26789 8375 26847 8381
rect 26881 8415 26939 8421
rect 26881 8381 26893 8415
rect 26927 8412 26939 8415
rect 27065 8415 27123 8421
rect 27065 8412 27077 8415
rect 26927 8384 27077 8412
rect 26927 8381 26939 8384
rect 26881 8375 26939 8381
rect 27065 8381 27077 8384
rect 27111 8381 27123 8415
rect 27065 8375 27123 8381
rect 27157 8415 27215 8421
rect 27157 8381 27169 8415
rect 27203 8412 27215 8415
rect 27341 8415 27399 8421
rect 27341 8412 27353 8415
rect 27203 8384 27353 8412
rect 27203 8381 27215 8384
rect 27157 8375 27215 8381
rect 27341 8381 27353 8384
rect 27387 8381 27399 8415
rect 27341 8375 27399 8381
rect 27433 8415 27491 8421
rect 27433 8381 27445 8415
rect 27479 8412 27491 8415
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 27479 8384 27629 8412
rect 27479 8381 27491 8384
rect 27433 8375 27491 8381
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 27709 8415 27767 8421
rect 27709 8381 27721 8415
rect 27755 8412 27767 8415
rect 27893 8415 27951 8421
rect 27893 8412 27905 8415
rect 27755 8384 27905 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 27893 8381 27905 8384
rect 27939 8381 27951 8415
rect 27893 8375 27951 8381
rect 27985 8415 28043 8421
rect 27985 8381 27997 8415
rect 28031 8412 28043 8415
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 28031 8384 28181 8412
rect 28031 8381 28043 8384
rect 27985 8375 28043 8381
rect 28169 8381 28181 8384
rect 28215 8381 28227 8415
rect 28169 8375 28227 8381
rect 28261 8415 28319 8421
rect 28261 8381 28273 8415
rect 28307 8412 28319 8415
rect 28445 8415 28503 8421
rect 28445 8412 28457 8415
rect 28307 8384 28457 8412
rect 28307 8381 28319 8384
rect 28261 8375 28319 8381
rect 28445 8381 28457 8384
rect 28491 8381 28503 8415
rect 28445 8375 28503 8381
rect 28537 8415 28595 8421
rect 28537 8381 28549 8415
rect 28583 8412 28595 8415
rect 28997 8415 29055 8421
rect 28997 8412 29009 8415
rect 28583 8384 29009 8412
rect 28583 8381 28595 8384
rect 28537 8375 28595 8381
rect 28997 8381 29009 8384
rect 29043 8381 29055 8415
rect 28997 8375 29055 8381
rect 24581 8347 24639 8353
rect 24581 8344 24593 8347
rect 24412 8316 24593 8344
rect 19291 8313 19303 8316
rect 19245 8307 19303 8313
rect 24581 8313 24593 8316
rect 24627 8313 24639 8347
rect 24581 8307 24639 8313
rect 26605 8347 26663 8353
rect 26605 8313 26617 8347
rect 26651 8344 26663 8347
rect 26804 8344 26832 8375
rect 29270 8372 29276 8424
rect 29328 8372 29334 8424
rect 26651 8316 26832 8344
rect 26651 8313 26663 8316
rect 26605 8307 26663 8313
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8276 7343 8279
rect 7466 8276 7472 8288
rect 7331 8248 7472 8276
rect 7331 8245 7343 8248
rect 7285 8239 7343 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7561 8279 7619 8285
rect 7561 8245 7573 8279
rect 7607 8276 7619 8279
rect 7742 8276 7748 8288
rect 7607 8248 7748 8276
rect 7607 8245 7619 8248
rect 7561 8239 7619 8245
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 8570 8236 8576 8288
rect 8628 8236 8634 8288
rect 8849 8279 8907 8285
rect 8849 8245 8861 8279
rect 8895 8276 8907 8279
rect 9030 8276 9036 8288
rect 8895 8248 9036 8276
rect 8895 8245 8907 8248
rect 8849 8239 8907 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 15436 8248 16037 8276
rect 15436 8236 15442 8248
rect 16025 8245 16037 8248
rect 16071 8245 16083 8279
rect 16025 8239 16083 8245
rect 29086 8236 29092 8288
rect 29144 8236 29150 8288
rect 552 8186 31648 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31648 8186
rect 552 8112 31648 8134
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8720 8044 9137 8072
rect 8720 8032 8726 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 17092 8044 17233 8072
rect 17092 8032 17098 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 24121 8075 24179 8081
rect 24121 8041 24133 8075
rect 24167 8072 24179 8075
rect 24486 8072 24492 8084
rect 24167 8044 24492 8072
rect 24167 8041 24179 8044
rect 24121 8035 24179 8041
rect 24486 8032 24492 8044
rect 24544 8032 24550 8084
rect 28721 8075 28779 8081
rect 28721 8041 28733 8075
rect 28767 8072 28779 8075
rect 29270 8072 29276 8084
rect 28767 8044 29276 8072
rect 28767 8041 28779 8044
rect 28721 8035 28779 8041
rect 29270 8032 29276 8044
rect 29328 8032 29334 8084
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 7432 7976 7849 8004
rect 7432 7964 7438 7976
rect 7837 7973 7849 7976
rect 7883 7973 7895 8007
rect 13725 8007 13783 8013
rect 13725 8004 13737 8007
rect 7837 7967 7895 7973
rect 13280 7976 13737 8004
rect 7466 7896 7472 7948
rect 7524 7896 7530 7948
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 8018 7896 8024 7948
rect 8076 7896 8082 7948
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 8159 7908 8309 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 8297 7905 8309 7908
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 8570 7896 8576 7948
rect 8628 7896 8634 7948
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 11238 7936 11244 7948
rect 10827 7908 11244 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 13280 7945 13308 7976
rect 13725 7973 13737 7976
rect 13771 7973 13783 8007
rect 16209 8007 16267 8013
rect 16209 8004 16221 8007
rect 13725 7967 13783 7973
rect 15120 7976 16221 8004
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11379 7908 11529 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11655 7908 11805 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11931 7908 12081 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12207 7908 12357 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12483 7908 12633 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12713 7939 12771 7945
rect 12713 7905 12725 7939
rect 12759 7936 12771 7939
rect 12897 7939 12955 7945
rect 12897 7936 12909 7939
rect 12759 7908 12909 7936
rect 12759 7905 12771 7908
rect 12713 7899 12771 7905
rect 12897 7905 12909 7908
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 13035 7908 13185 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13538 7896 13544 7948
rect 13596 7896 13602 7948
rect 15120 7945 15148 7976
rect 16209 7973 16221 7976
rect 16255 7973 16267 8007
rect 16209 7967 16267 7973
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 8536 7840 8677 7868
rect 8536 7828 8542 7840
rect 8665 7837 8677 7840
rect 8711 7837 8723 7871
rect 8665 7831 8723 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13648 7868 13676 7899
rect 15378 7896 15384 7948
rect 15436 7896 15442 7948
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7905 15531 7939
rect 15473 7899 15531 7905
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15611 7908 15761 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 15887 7908 16129 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7936 17371 7939
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 17359 7908 17509 7936
rect 17359 7905 17371 7908
rect 17313 7899 17371 7905
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17773 7939 17831 7945
rect 17773 7936 17785 7939
rect 17635 7908 17785 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17773 7905 17785 7908
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 17911 7908 18061 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 18187 7908 18337 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7936 18475 7939
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 18463 7908 18613 7936
rect 18463 7905 18475 7908
rect 18417 7899 18475 7905
rect 18601 7905 18613 7908
rect 18647 7905 18659 7939
rect 18601 7899 18659 7905
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 18739 7908 18889 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 13495 7840 13676 7868
rect 15289 7871 15347 7877
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15488 7868 15516 7899
rect 18966 7896 18972 7948
rect 19024 7896 19030 7948
rect 20346 7896 20352 7948
rect 20404 7896 20410 7948
rect 20441 7939 20499 7945
rect 20441 7905 20453 7939
rect 20487 7905 20499 7939
rect 20441 7899 20499 7905
rect 20533 7939 20591 7945
rect 20533 7905 20545 7939
rect 20579 7936 20591 7939
rect 20717 7939 20775 7945
rect 20717 7936 20729 7939
rect 20579 7908 20729 7936
rect 20579 7905 20591 7908
rect 20533 7899 20591 7905
rect 20717 7905 20729 7908
rect 20763 7905 20775 7939
rect 20717 7899 20775 7905
rect 20809 7939 20867 7945
rect 20809 7905 20821 7939
rect 20855 7936 20867 7939
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 20855 7908 21281 7936
rect 20855 7905 20867 7908
rect 20809 7899 20867 7905
rect 21269 7905 21281 7908
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 21361 7939 21419 7945
rect 21361 7905 21373 7939
rect 21407 7936 21419 7939
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 21407 7908 21557 7936
rect 21407 7905 21419 7908
rect 21361 7899 21419 7905
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21637 7939 21695 7945
rect 21637 7905 21649 7939
rect 21683 7936 21695 7939
rect 21821 7939 21879 7945
rect 21821 7936 21833 7939
rect 21683 7908 21833 7936
rect 21683 7905 21695 7908
rect 21637 7899 21695 7905
rect 21821 7905 21833 7908
rect 21867 7905 21879 7939
rect 21821 7899 21879 7905
rect 21913 7939 21971 7945
rect 21913 7905 21925 7939
rect 21959 7936 21971 7939
rect 22097 7939 22155 7945
rect 22097 7936 22109 7939
rect 21959 7908 22109 7936
rect 21959 7905 21971 7908
rect 21913 7899 21971 7905
rect 22097 7905 22109 7908
rect 22143 7905 22155 7939
rect 22097 7899 22155 7905
rect 22189 7939 22247 7945
rect 22189 7905 22201 7939
rect 22235 7936 22247 7939
rect 22373 7939 22431 7945
rect 22373 7936 22385 7939
rect 22235 7908 22385 7936
rect 22235 7905 22247 7908
rect 22189 7899 22247 7905
rect 22373 7905 22385 7908
rect 22419 7905 22431 7939
rect 22373 7899 22431 7905
rect 15335 7840 15516 7868
rect 20257 7871 20315 7877
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20456 7868 20484 7899
rect 22646 7896 22652 7948
rect 22704 7896 22710 7948
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 22925 7939 22983 7945
rect 22925 7936 22937 7939
rect 22787 7908 22937 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 22925 7905 22937 7908
rect 22971 7905 22983 7939
rect 22925 7899 22983 7905
rect 23017 7939 23075 7945
rect 23017 7905 23029 7939
rect 23063 7936 23075 7939
rect 23201 7939 23259 7945
rect 23201 7936 23213 7939
rect 23063 7908 23213 7936
rect 23063 7905 23075 7908
rect 23017 7899 23075 7905
rect 23201 7905 23213 7908
rect 23247 7905 23259 7939
rect 23201 7899 23259 7905
rect 23474 7896 23480 7948
rect 23532 7896 23538 7948
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7936 24271 7939
rect 24397 7939 24455 7945
rect 24397 7936 24409 7939
rect 24259 7908 24409 7936
rect 24259 7905 24271 7908
rect 24213 7899 24271 7905
rect 24397 7905 24409 7908
rect 24443 7905 24455 7939
rect 24397 7899 24455 7905
rect 24489 7939 24547 7945
rect 24489 7905 24501 7939
rect 24535 7936 24547 7939
rect 24673 7939 24731 7945
rect 24673 7936 24685 7939
rect 24535 7908 24685 7936
rect 24535 7905 24547 7908
rect 24489 7899 24547 7905
rect 24673 7905 24685 7908
rect 24719 7905 24731 7939
rect 24673 7899 24731 7905
rect 24765 7939 24823 7945
rect 24765 7905 24777 7939
rect 24811 7936 24823 7939
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24811 7908 24961 7936
rect 24811 7905 24823 7908
rect 24765 7899 24823 7905
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 25041 7939 25099 7945
rect 25041 7905 25053 7939
rect 25087 7936 25099 7939
rect 25225 7939 25283 7945
rect 25225 7936 25237 7939
rect 25087 7908 25237 7936
rect 25087 7905 25099 7908
rect 25041 7899 25099 7905
rect 25225 7905 25237 7908
rect 25271 7905 25283 7939
rect 25225 7899 25283 7905
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7936 25375 7939
rect 25501 7939 25559 7945
rect 25501 7936 25513 7939
rect 25363 7908 25513 7936
rect 25363 7905 25375 7908
rect 25317 7899 25375 7905
rect 25501 7905 25513 7908
rect 25547 7905 25559 7939
rect 25501 7899 25559 7905
rect 25593 7939 25651 7945
rect 25593 7905 25605 7939
rect 25639 7936 25651 7939
rect 25777 7939 25835 7945
rect 25777 7936 25789 7939
rect 25639 7908 25789 7936
rect 25639 7905 25651 7908
rect 25593 7899 25651 7905
rect 25777 7905 25789 7908
rect 25823 7905 25835 7939
rect 25777 7899 25835 7905
rect 25869 7939 25927 7945
rect 25869 7905 25881 7939
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 20303 7840 20484 7868
rect 25884 7868 25912 7899
rect 25958 7896 25964 7948
rect 26016 7896 26022 7948
rect 28813 7939 28871 7945
rect 28813 7905 28825 7939
rect 28859 7936 28871 7939
rect 28997 7939 29055 7945
rect 28997 7936 29009 7939
rect 28859 7908 29009 7936
rect 28859 7905 28871 7908
rect 28813 7899 28871 7905
rect 28997 7905 29009 7908
rect 29043 7905 29055 7939
rect 28997 7899 29055 7905
rect 29086 7896 29092 7948
rect 29144 7896 29150 7948
rect 26053 7871 26111 7877
rect 26053 7868 26065 7871
rect 25884 7840 26065 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 26053 7837 26065 7840
rect 26099 7837 26111 7871
rect 26053 7831 26111 7837
rect 23014 7760 23020 7812
rect 23072 7800 23078 7812
rect 23569 7803 23627 7809
rect 23569 7800 23581 7803
rect 23072 7772 23581 7800
rect 23072 7760 23078 7772
rect 23569 7769 23581 7772
rect 23615 7769 23627 7803
rect 23569 7763 23627 7769
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 7432 7704 8401 7732
rect 7432 7692 7438 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 8389 7695 8447 7701
rect 11241 7735 11299 7741
rect 11241 7701 11253 7735
rect 11287 7732 11299 7735
rect 11330 7732 11336 7744
rect 11287 7704 11336 7732
rect 11287 7701 11299 7704
rect 11241 7695 11299 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 15013 7735 15071 7741
rect 15013 7701 15025 7735
rect 15059 7732 15071 7735
rect 15194 7732 15200 7744
rect 15059 7704 15200 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 22465 7735 22523 7741
rect 22465 7732 22477 7735
rect 21968 7704 22477 7732
rect 21968 7692 21974 7704
rect 22465 7701 22477 7704
rect 22511 7701 22523 7735
rect 22465 7695 22523 7701
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 23293 7735 23351 7741
rect 23293 7732 23305 7735
rect 22796 7704 23305 7732
rect 22796 7692 22802 7704
rect 23293 7701 23305 7704
rect 23339 7701 23351 7735
rect 23293 7695 23351 7701
rect 552 7642 31648 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31648 7642
rect 552 7568 31648 7590
rect 11238 7488 11244 7540
rect 11296 7488 11302 7540
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13596 7500 13645 7528
rect 13596 7488 13602 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 20533 7531 20591 7537
rect 20533 7528 20545 7531
rect 20404 7500 20545 7528
rect 20404 7488 20410 7500
rect 20533 7497 20545 7500
rect 20579 7497 20591 7531
rect 20533 7491 20591 7497
rect 21821 7531 21879 7537
rect 21821 7497 21833 7531
rect 21867 7528 21879 7531
rect 22646 7528 22652 7540
rect 21867 7500 22652 7528
rect 21867 7497 21879 7500
rect 21821 7491 21879 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 25317 7531 25375 7537
rect 25317 7497 25329 7531
rect 25363 7528 25375 7531
rect 25958 7528 25964 7540
rect 25363 7500 25964 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7429 17279 7463
rect 17221 7423 17279 7429
rect 19981 7463 20039 7469
rect 19981 7429 19993 7463
rect 20027 7460 20039 7463
rect 23474 7460 23480 7472
rect 20027 7432 20484 7460
rect 20027 7429 20039 7432
rect 19981 7423 20039 7429
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 9585 7395 9643 7401
rect 7607 7364 7788 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7147 7296 7297 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7374 7284 7380 7336
rect 7432 7284 7438 7336
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7760 7333 7788 7364
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 9631 7364 10088 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 10060 7333 10088 7364
rect 11348 7364 11529 7392
rect 11348 7333 11376 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 11517 7355 11575 7361
rect 14016 7364 14197 7392
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7883 7296 8033 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8159 7296 8401 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 8527 7296 8677 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8803 7296 8953 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9079 7296 9229 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 9355 7296 9505 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 11333 7327 11391 7333
rect 11333 7293 11345 7327
rect 11379 7293 11391 7327
rect 11333 7287 11391 7293
rect 9968 7256 9996 7287
rect 11422 7284 11428 7336
rect 11480 7284 11486 7336
rect 14016 7333 14044 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 17236 7392 17264 7423
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 17236 7364 17448 7392
rect 14185 7355 14243 7361
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13771 7296 13921 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14090 7284 14096 7336
rect 14148 7284 14154 7336
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15335 7296 15485 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15611 7296 15761 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 17218 7324 17224 7336
rect 17175 7296 17224 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 17420 7333 17448 7364
rect 20088 7364 20269 7392
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 17543 7296 17693 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 19794 7284 19800 7336
rect 19852 7284 19858 7336
rect 20088 7333 20116 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20456 7333 20484 7432
rect 22664 7432 23480 7460
rect 22664 7401 22692 7432
rect 23474 7420 23480 7432
rect 23532 7420 23538 7472
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 25869 7395 25927 7401
rect 25869 7392 25881 7395
rect 22971 7364 23152 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9968 7228 10149 7256
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 19705 7259 19763 7265
rect 19705 7225 19717 7259
rect 19751 7256 19763 7259
rect 20180 7256 20208 7287
rect 21910 7284 21916 7336
rect 21968 7284 21974 7336
rect 22738 7284 22744 7336
rect 22796 7284 22802 7336
rect 23014 7284 23020 7336
rect 23072 7284 23078 7336
rect 23124 7333 23152 7364
rect 25700 7364 25881 7392
rect 25700 7333 25728 7364
rect 25869 7361 25881 7364
rect 25915 7361 25927 7395
rect 25869 7355 25927 7361
rect 23109 7327 23167 7333
rect 23109 7293 23121 7327
rect 23155 7293 23167 7327
rect 23109 7287 23167 7293
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7324 23259 7327
rect 23385 7327 23443 7333
rect 23385 7324 23397 7327
rect 23247 7296 23397 7324
rect 23247 7293 23259 7296
rect 23201 7287 23259 7293
rect 23385 7293 23397 7296
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 25409 7327 25467 7333
rect 25409 7293 25421 7327
rect 25455 7324 25467 7327
rect 25593 7327 25651 7333
rect 25593 7324 25605 7327
rect 25455 7296 25605 7324
rect 25455 7293 25467 7296
rect 25409 7287 25467 7293
rect 25593 7293 25605 7296
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 25685 7327 25743 7333
rect 25685 7293 25697 7327
rect 25731 7293 25743 7327
rect 25685 7287 25743 7293
rect 25774 7284 25780 7336
rect 25832 7284 25838 7336
rect 19751 7228 20208 7256
rect 19751 7225 19763 7228
rect 19705 7219 19763 7225
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7742 7188 7748 7200
rect 7055 7160 7748 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 9950 7188 9956 7200
rect 9907 7160 9956 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15252 7160 15853 7188
rect 15252 7148 15258 7160
rect 15841 7157 15853 7160
rect 15887 7157 15899 7191
rect 15841 7151 15899 7157
rect 17770 7148 17776 7200
rect 17828 7148 17834 7200
rect 18141 7191 18199 7197
rect 18141 7157 18153 7191
rect 18187 7188 18199 7191
rect 18230 7188 18236 7200
rect 18187 7160 18236 7188
rect 18187 7157 18199 7160
rect 18141 7151 18199 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 23474 7148 23480 7200
rect 23532 7148 23538 7200
rect 552 7098 31648 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31648 7098
rect 552 7024 31648 7046
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7708 6956 7849 6984
rect 7708 6944 7714 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 17129 6987 17187 6993
rect 17129 6953 17141 6987
rect 17175 6984 17187 6987
rect 17218 6984 17224 6996
rect 17175 6956 17224 6984
rect 17175 6953 17187 6956
rect 17129 6947 17187 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 19794 6944 19800 6996
rect 19852 6944 19858 6996
rect 25317 6987 25375 6993
rect 25317 6953 25329 6987
rect 25363 6984 25375 6987
rect 25774 6984 25780 6996
rect 25363 6956 25780 6984
rect 25363 6953 25375 6956
rect 25317 6947 25375 6953
rect 25774 6944 25780 6956
rect 25832 6944 25838 6996
rect 23474 6916 23480 6928
rect 16684 6888 17172 6916
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6687 6820 6837 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6963 6820 7113 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 7742 6808 7748 6860
rect 7800 6808 7806 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 9876 6780 9904 6811
rect 9950 6808 9956 6860
rect 10008 6808 10014 6860
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 10091 6820 10241 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10367 6820 10517 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 13446 6808 13452 6860
rect 13504 6808 13510 6860
rect 13725 6851 13783 6857
rect 13725 6817 13737 6851
rect 13771 6848 13783 6851
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13771 6820 13921 6848
rect 13771 6817 13783 6820
rect 13725 6811 13783 6817
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 13909 6811 13967 6817
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6848 14059 6851
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14047 6820 14197 6848
rect 14047 6817 14059 6820
rect 14001 6811 14059 6817
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 14277 6851 14335 6857
rect 14277 6817 14289 6851
rect 14323 6848 14335 6851
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14323 6820 14473 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14599 6820 14749 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 9876 6752 10609 6780
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 14090 6780 14096 6792
rect 13403 6752 14096 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14844 6712 14872 6811
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15304 6780 15332 6811
rect 15930 6808 15936 6860
rect 15988 6808 15994 6860
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16347 6820 16497 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 16684 6848 16712 6888
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16623 6820 16712 6848
rect 16776 6820 16957 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 15151 6752 15332 6780
rect 15841 6783 15899 6789
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 16224 6780 16252 6811
rect 15887 6752 16252 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 15381 6715 15439 6721
rect 15381 6712 15393 6715
rect 14844 6684 15393 6712
rect 15381 6681 15393 6684
rect 15427 6681 15439 6715
rect 16776 6712 16804 6820
rect 16945 6817 16957 6820
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 17037 6851 17095 6857
rect 17037 6817 17049 6851
rect 17083 6817 17095 6851
rect 17144 6848 17172 6888
rect 19812 6888 20024 6916
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 17144 6820 17325 6848
rect 17037 6811 17095 6817
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6780 16911 6783
rect 17052 6780 17080 6811
rect 17770 6808 17776 6860
rect 17828 6808 17834 6860
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 18046 6848 18052 6860
rect 17911 6820 18052 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18325 6851 18383 6857
rect 18325 6817 18337 6851
rect 18371 6848 18383 6851
rect 18601 6851 18659 6857
rect 18601 6848 18613 6851
rect 18371 6820 18613 6848
rect 18371 6817 18383 6820
rect 18325 6811 18383 6817
rect 18601 6817 18613 6820
rect 18647 6817 18659 6851
rect 18601 6811 18659 6817
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6848 18751 6851
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18739 6820 18889 6848
rect 18739 6817 18751 6820
rect 18693 6811 18751 6817
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 18969 6851 19027 6857
rect 18969 6817 18981 6851
rect 19015 6848 19027 6851
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 19015 6820 19165 6848
rect 19015 6817 19027 6820
rect 18969 6811 19027 6817
rect 19153 6817 19165 6820
rect 19199 6817 19211 6851
rect 19153 6811 19211 6817
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 19291 6820 19441 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6848 19579 6851
rect 19812 6848 19840 6888
rect 19996 6857 20024 6888
rect 23124 6888 23480 6916
rect 23124 6857 23152 6888
rect 23474 6876 23480 6888
rect 23532 6876 23538 6928
rect 19567 6820 19840 6848
rect 19889 6851 19947 6857
rect 19567 6817 19579 6820
rect 19521 6811 19579 6817
rect 19889 6817 19901 6851
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 22051 6820 22201 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22189 6817 22201 6820
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 22281 6851 22339 6857
rect 22281 6817 22293 6851
rect 22327 6848 22339 6851
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 22327 6820 22477 6848
rect 22327 6817 22339 6820
rect 22281 6811 22339 6817
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6848 22615 6851
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22603 6820 22753 6848
rect 22603 6817 22615 6820
rect 22557 6811 22615 6817
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 22741 6811 22799 6817
rect 22833 6851 22891 6857
rect 22833 6817 22845 6851
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6817 23167 6851
rect 23109 6811 23167 6817
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6817 23259 6851
rect 23201 6811 23259 6817
rect 25409 6851 25467 6857
rect 25409 6817 25421 6851
rect 25455 6848 25467 6851
rect 25593 6851 25651 6857
rect 25593 6848 25605 6851
rect 25455 6820 25605 6848
rect 25455 6817 25467 6820
rect 25409 6811 25467 6817
rect 25593 6817 25605 6820
rect 25639 6817 25651 6851
rect 25593 6811 25651 6817
rect 25685 6851 25743 6857
rect 25685 6817 25697 6851
rect 25731 6848 25743 6851
rect 25869 6851 25927 6857
rect 25869 6848 25881 6851
rect 25731 6820 25881 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 25869 6817 25881 6820
rect 25915 6817 25927 6851
rect 25869 6811 25927 6817
rect 25961 6851 26019 6857
rect 25961 6817 25973 6851
rect 26007 6817 26019 6851
rect 25961 6811 26019 6817
rect 16899 6752 17080 6780
rect 19904 6780 19932 6811
rect 20073 6783 20131 6789
rect 20073 6780 20085 6783
rect 19904 6752 20085 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 20073 6749 20085 6752
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 16776 6684 17417 6712
rect 15381 6675 15439 6681
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 22848 6712 22876 6811
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6780 23075 6783
rect 23216 6780 23244 6811
rect 23063 6752 23244 6780
rect 25976 6780 26004 6811
rect 26050 6808 26056 6860
rect 26108 6808 26114 6860
rect 26145 6783 26203 6789
rect 26145 6780 26157 6783
rect 25976 6752 26157 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 26145 6749 26157 6752
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 23293 6715 23351 6721
rect 23293 6712 23305 6715
rect 22848 6684 23305 6712
rect 17405 6675 17463 6681
rect 23293 6681 23305 6684
rect 23339 6681 23351 6715
rect 23293 6675 23351 6681
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 6512 6616 6561 6644
rect 6512 6604 6518 6616
rect 6549 6613 6561 6616
rect 6595 6613 6607 6647
rect 6549 6607 6607 6613
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10042 6644 10048 6656
rect 9815 6616 10048 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 13630 6604 13636 6656
rect 13688 6604 13694 6656
rect 21910 6604 21916 6656
rect 21968 6604 21974 6656
rect 552 6554 31648 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31648 6554
rect 552 6480 31648 6502
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13504 6412 13737 6440
rect 13504 6400 13510 6412
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15988 6412 16221 6440
rect 15988 6400 15994 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16209 6403 16267 6409
rect 25317 6443 25375 6449
rect 25317 6409 25329 6443
rect 25363 6440 25375 6443
rect 26050 6440 26056 6452
rect 25363 6412 26056 6440
rect 25363 6409 25375 6412
rect 25317 6403 25375 6409
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 21545 6375 21603 6381
rect 21545 6341 21557 6375
rect 21591 6372 21603 6375
rect 21591 6344 22600 6372
rect 21591 6341 21603 6344
rect 21545 6335 21603 6341
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 5920 6276 6653 6304
rect 5920 6245 5948 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 6641 6267 6699 6273
rect 8128 6276 8493 6304
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 6227 6208 6377 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6454 6196 6460 6248
rect 6512 6196 6518 6248
rect 8128 6245 8156 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 11655 6276 11836 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 7331 6208 7481 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 7469 6205 7481 6208
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6236 7619 6239
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7607 6208 7757 6236
rect 7607 6205 7619 6208
rect 7561 6199 7619 6205
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7883 6208 8033 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 6089 6171 6147 6177
rect 6089 6137 6101 6171
rect 6135 6168 6147 6171
rect 6564 6168 6592 6199
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 8260 6208 8401 6236
rect 8260 6196 8266 6208
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10321 6239 10379 6245
rect 10321 6236 10333 6239
rect 10183 6208 10333 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 10321 6205 10333 6208
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 11146 6196 11152 6248
rect 11204 6196 11210 6248
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 6135 6140 6592 6168
rect 11057 6171 11115 6177
rect 6135 6137 6147 6140
rect 6089 6131 6147 6137
rect 11057 6137 11069 6171
rect 11103 6168 11115 6171
rect 11256 6168 11284 6199
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 11808 6245 11836 6276
rect 12912 6276 13093 6304
rect 12912 6245 12940 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 13081 6267 13139 6273
rect 16316 6276 16497 6304
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11931 6208 12081 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 12207 6208 12357 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 11103 6140 11284 6168
rect 12437 6171 12495 6177
rect 11103 6137 11115 6140
rect 11057 6131 11115 6137
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 13004 6168 13032 6199
rect 13630 6196 13636 6248
rect 13688 6196 13694 6248
rect 16316 6245 16344 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 22373 6307 22431 6313
rect 22373 6304 22385 6307
rect 16485 6267 16543 6273
rect 21652 6276 22385 6304
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15856 6208 16037 6236
rect 12483 6140 13032 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 10284 6072 10425 6100
rect 10284 6060 10290 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11790 6100 11796 6112
rect 11379 6072 11796 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12676 6072 12817 6100
rect 12676 6060 12682 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 15856 6100 15884 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 15933 6171 15991 6177
rect 15933 6137 15945 6171
rect 15979 6168 15991 6171
rect 16408 6168 16436 6199
rect 16666 6196 16672 6248
rect 16724 6196 16730 6248
rect 21652 6245 21680 6276
rect 22373 6273 22385 6276
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 21637 6239 21695 6245
rect 21637 6205 21649 6239
rect 21683 6205 21695 6239
rect 21637 6199 21695 6205
rect 21910 6196 21916 6248
rect 21968 6196 21974 6248
rect 22572 6245 22600 6344
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6205 22063 6239
rect 22005 6199 22063 6205
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22281 6239 22339 6245
rect 22281 6236 22293 6239
rect 22143 6208 22293 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22281 6205 22293 6208
rect 22327 6205 22339 6239
rect 22281 6199 22339 6205
rect 22557 6239 22615 6245
rect 22557 6205 22569 6239
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 25409 6239 25467 6245
rect 25409 6205 25421 6239
rect 25455 6236 25467 6239
rect 25593 6239 25651 6245
rect 25593 6236 25605 6239
rect 25455 6208 25605 6236
rect 25455 6205 25467 6208
rect 25409 6199 25467 6205
rect 25593 6205 25605 6208
rect 25639 6205 25651 6239
rect 25593 6199 25651 6205
rect 25685 6239 25743 6245
rect 25685 6205 25697 6239
rect 25731 6236 25743 6239
rect 25869 6239 25927 6245
rect 25869 6236 25881 6239
rect 25731 6208 25881 6236
rect 25731 6205 25743 6208
rect 25685 6199 25743 6205
rect 25869 6205 25881 6208
rect 25915 6205 25927 6239
rect 25869 6199 25927 6205
rect 25961 6239 26019 6245
rect 25961 6205 25973 6239
rect 26007 6205 26019 6239
rect 25961 6199 26019 6205
rect 15979 6140 16436 6168
rect 21821 6171 21879 6177
rect 15979 6137 15991 6140
rect 15933 6131 15991 6137
rect 21821 6137 21833 6171
rect 21867 6168 21879 6171
rect 22020 6168 22048 6199
rect 21867 6140 22048 6168
rect 25976 6168 26004 6199
rect 26050 6196 26056 6248
rect 26108 6196 26114 6248
rect 26145 6171 26203 6177
rect 26145 6168 26157 6171
rect 25976 6140 26157 6168
rect 21867 6137 21879 6140
rect 21821 6131 21879 6137
rect 26145 6137 26157 6140
rect 26191 6137 26203 6171
rect 26145 6131 26203 6137
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 15856 6072 16773 6100
rect 12805 6063 12863 6069
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 16761 6063 16819 6069
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22060 6072 22661 6100
rect 22060 6060 22066 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 552 6010 31648 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31648 6010
rect 552 5936 31648 5958
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11333 5899 11391 5905
rect 11333 5896 11345 5899
rect 11204 5868 11345 5896
rect 11204 5856 11210 5868
rect 11333 5865 11345 5868
rect 11379 5865 11391 5899
rect 11333 5859 11391 5865
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11756 5868 11897 5896
rect 11756 5856 11762 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16666 5896 16672 5908
rect 15887 5868 16672 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 25317 5899 25375 5905
rect 25317 5865 25329 5899
rect 25363 5896 25375 5899
rect 26050 5896 26056 5908
rect 25363 5868 26056 5896
rect 25363 5865 25375 5868
rect 25317 5859 25375 5865
rect 26050 5856 26056 5868
rect 26108 5856 26114 5908
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6472 5800 6653 5828
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 5644 5692 5672 5723
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 6472 5769 6500 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 9585 5831 9643 5837
rect 9585 5828 9597 5831
rect 6641 5791 6699 5797
rect 9140 5800 9597 5828
rect 9140 5769 9168 5800
rect 9585 5797 9597 5800
rect 9631 5797 9643 5831
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 9585 5791 9643 5797
rect 11164 5800 11621 5828
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8343 5732 8493 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 8481 5723 8539 5729
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 8849 5763 8907 5769
rect 8849 5729 8861 5763
rect 8895 5760 8907 5763
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8895 5732 9045 5760
rect 8895 5729 8907 5732
rect 8849 5723 8907 5729
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5644 5664 5917 5692
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 5537 5627 5595 5633
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 6564 5624 6592 5723
rect 5583 5596 6592 5624
rect 8588 5624 8616 5723
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 9232 5692 9260 5723
rect 9490 5720 9496 5772
rect 9548 5720 9554 5772
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 9999 5732 10149 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10226 5720 10232 5772
rect 10284 5720 10290 5772
rect 11164 5769 11192 5800
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11609 5791 11667 5797
rect 12529 5831 12587 5837
rect 12529 5797 12541 5831
rect 12575 5828 12587 5831
rect 13909 5831 13967 5837
rect 12575 5800 12756 5828
rect 12575 5797 12587 5800
rect 12529 5791 12587 5797
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 10459 5732 10609 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10597 5729 10609 5732
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11241 5723 11299 5729
rect 11348 5732 11529 5760
rect 8803 5664 9260 5692
rect 9861 5695 9919 5701
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 10336 5692 10364 5723
rect 9907 5664 10364 5692
rect 11057 5695 11115 5701
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11256 5692 11284 5723
rect 11103 5664 11284 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8588 5596 9321 5624
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 10689 5627 10747 5633
rect 10689 5593 10701 5627
rect 10735 5624 10747 5627
rect 11348 5624 11376 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11790 5720 11796 5772
rect 11848 5720 11854 5772
rect 12618 5720 12624 5772
rect 12676 5720 12682 5772
rect 12728 5769 12756 5800
rect 13909 5797 13921 5831
rect 13955 5828 13967 5831
rect 16485 5831 16543 5837
rect 16485 5828 16497 5831
rect 13955 5800 14504 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 14476 5769 14504 5800
rect 16316 5800 16497 5828
rect 16316 5769 16344 5800
rect 16485 5797 16497 5800
rect 16531 5797 16543 5831
rect 25869 5831 25927 5837
rect 25869 5828 25881 5831
rect 16485 5791 16543 5797
rect 25700 5800 25881 5828
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12851 5732 13001 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 13127 5732 13277 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13403 5732 13553 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5760 13691 5763
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 13679 5732 13829 5760
rect 13679 5729 13691 5732
rect 13633 5723 13691 5729
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 15979 5732 16221 5760
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 14384 5692 14412 5723
rect 16390 5720 16396 5772
rect 16448 5720 16454 5772
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 17359 5732 17509 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5760 17647 5763
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17635 5732 17785 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 17773 5729 17785 5732
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 17911 5732 18061 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18049 5723 18107 5729
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5760 18199 5763
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18187 5732 18337 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5760 18475 5763
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18463 5732 18613 5760
rect 18463 5729 18475 5732
rect 18417 5723 18475 5729
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 18877 5763 18935 5769
rect 18877 5760 18889 5763
rect 18739 5732 18889 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 18877 5729 18889 5732
rect 18923 5729 18935 5763
rect 18877 5723 18935 5729
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5760 19027 5763
rect 19153 5763 19211 5769
rect 19153 5760 19165 5763
rect 19015 5732 19165 5760
rect 19015 5729 19027 5732
rect 18969 5723 19027 5729
rect 19153 5729 19165 5732
rect 19199 5729 19211 5763
rect 19153 5723 19211 5729
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19337 5763 19395 5769
rect 19337 5729 19349 5763
rect 19383 5760 19395 5763
rect 19610 5760 19616 5772
rect 19383 5732 19616 5760
rect 19383 5729 19395 5732
rect 19337 5723 19395 5729
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14384 5664 14565 5692
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 19260 5692 19288 5723
rect 19610 5720 19616 5732
rect 19668 5720 19674 5772
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 19981 5763 20039 5769
rect 19981 5760 19993 5763
rect 19843 5732 19993 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 19981 5729 19993 5732
rect 20027 5729 20039 5763
rect 19981 5723 20039 5729
rect 20073 5763 20131 5769
rect 20073 5729 20085 5763
rect 20119 5760 20131 5763
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 20119 5732 20269 5760
rect 20119 5729 20131 5732
rect 20073 5723 20131 5729
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 20349 5763 20407 5769
rect 20349 5729 20361 5763
rect 20395 5729 20407 5763
rect 20349 5723 20407 5729
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19260 5664 19441 5692
rect 14553 5655 14611 5661
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 20364 5692 20392 5723
rect 20438 5720 20444 5772
rect 20496 5720 20502 5772
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5760 20775 5763
rect 20806 5760 20812 5772
rect 20763 5732 20812 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 22002 5720 22008 5772
rect 22060 5720 22066 5772
rect 22097 5763 22155 5769
rect 22097 5729 22109 5763
rect 22143 5729 22155 5763
rect 22097 5723 22155 5729
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5760 22247 5763
rect 22373 5763 22431 5769
rect 22373 5760 22385 5763
rect 22235 5732 22385 5760
rect 22235 5729 22247 5732
rect 22189 5723 22247 5729
rect 22373 5729 22385 5732
rect 22419 5729 22431 5763
rect 22373 5723 22431 5729
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22511 5732 22661 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 22649 5723 22707 5729
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 20364 5664 20545 5692
rect 19429 5655 19487 5661
rect 20533 5661 20545 5664
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5692 21971 5695
rect 22112 5692 22140 5723
rect 24946 5720 24952 5772
rect 25004 5720 25010 5772
rect 25700 5769 25728 5800
rect 25869 5797 25881 5800
rect 25915 5797 25927 5831
rect 25869 5791 25927 5797
rect 25409 5763 25467 5769
rect 25409 5729 25421 5763
rect 25455 5760 25467 5763
rect 25593 5763 25651 5769
rect 25593 5760 25605 5763
rect 25455 5732 25605 5760
rect 25455 5729 25467 5732
rect 25409 5723 25467 5729
rect 25593 5729 25605 5732
rect 25639 5729 25651 5763
rect 25593 5723 25651 5729
rect 25685 5763 25743 5769
rect 25685 5729 25697 5763
rect 25731 5729 25743 5763
rect 25685 5723 25743 5729
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5729 25835 5763
rect 25777 5723 25835 5729
rect 21959 5664 22140 5692
rect 25041 5695 25099 5701
rect 21959 5661 21971 5664
rect 21913 5655 21971 5661
rect 25041 5661 25053 5695
rect 25087 5692 25099 5695
rect 25792 5692 25820 5723
rect 25087 5664 25820 5692
rect 25087 5661 25099 5664
rect 25041 5655 25099 5661
rect 10735 5596 11376 5624
rect 10735 5593 10747 5596
rect 10689 5587 10747 5593
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6454 5556 6460 5568
rect 6411 5528 6460 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 14274 5516 14280 5568
rect 14332 5516 14338 5568
rect 17126 5516 17132 5568
rect 17184 5556 17190 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 17184 5528 17233 5556
rect 17184 5516 17190 5528
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 17221 5519 17279 5525
rect 19702 5516 19708 5568
rect 19760 5516 19766 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 20809 5559 20867 5565
rect 20809 5556 20821 5559
rect 20772 5528 20821 5556
rect 20772 5516 20778 5528
rect 20809 5525 20821 5528
rect 20855 5525 20867 5559
rect 20809 5519 20867 5525
rect 22462 5516 22468 5568
rect 22520 5556 22526 5568
rect 22741 5559 22799 5565
rect 22741 5556 22753 5559
rect 22520 5528 22753 5556
rect 22520 5516 22526 5528
rect 22741 5525 22753 5528
rect 22787 5525 22799 5559
rect 22741 5519 22799 5525
rect 552 5466 31648 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31648 5466
rect 552 5392 31648 5414
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 9490 5352 9496 5364
rect 9079 5324 9496 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 15933 5355 15991 5361
rect 15933 5321 15945 5355
rect 15979 5352 15991 5355
rect 16390 5352 16396 5364
rect 15979 5324 16396 5352
rect 15979 5321 15991 5324
rect 15933 5315 15991 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 18785 5355 18843 5361
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 19610 5352 19616 5364
rect 18831 5324 19616 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 20257 5355 20315 5361
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 20806 5352 20812 5364
rect 20303 5324 20812 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5284 6883 5287
rect 14369 5287 14427 5293
rect 6871 5256 7328 5284
rect 6871 5253 6883 5256
rect 6825 5247 6883 5253
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6932 5188 7113 5216
rect 6454 5108 6460 5160
rect 6512 5108 6518 5160
rect 6932 5157 6960 5188
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 7300 5157 7328 5256
rect 14369 5253 14381 5287
rect 14415 5284 14427 5287
rect 19889 5287 19947 5293
rect 14415 5256 15148 5284
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 14752 5188 14964 5216
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9171 5120 9321 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 6549 5083 6607 5089
rect 6549 5049 6561 5083
rect 6595 5080 6607 5083
rect 7024 5080 7052 5111
rect 6595 5052 7052 5080
rect 9416 5080 9444 5111
rect 9490 5108 9496 5160
rect 9548 5108 9554 5160
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 14752 5157 14780 5188
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 9585 5083 9643 5089
rect 9585 5080 9597 5083
rect 9416 5052 9597 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 9585 5049 9597 5052
rect 9631 5049 9643 5083
rect 9585 5043 9643 5049
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 14844 5080 14872 5111
rect 14691 5052 14872 5080
rect 14936 5080 14964 5188
rect 15120 5157 15148 5256
rect 19889 5253 19901 5287
rect 19935 5284 19947 5287
rect 20438 5284 20444 5296
rect 19935 5256 20444 5284
rect 19935 5253 19947 5256
rect 19889 5247 19947 5253
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 20714 5216 20720 5228
rect 19996 5188 20720 5216
rect 15105 5151 15163 5157
rect 15105 5117 15117 5151
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 16025 5151 16083 5157
rect 16025 5117 16037 5151
rect 16071 5148 16083 5151
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 16071 5120 16221 5148
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 16209 5117 16221 5120
rect 16255 5117 16267 5151
rect 16209 5111 16267 5117
rect 16301 5151 16359 5157
rect 16301 5117 16313 5151
rect 16347 5148 16359 5151
rect 16485 5151 16543 5157
rect 16485 5148 16497 5151
rect 16347 5120 16497 5148
rect 16347 5117 16359 5120
rect 16301 5111 16359 5117
rect 16485 5117 16497 5120
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5148 16635 5151
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16623 5120 16773 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17037 5151 17095 5157
rect 17037 5148 17049 5151
rect 16899 5120 17049 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17037 5117 17049 5120
rect 17083 5117 17095 5151
rect 17037 5111 17095 5117
rect 17126 5108 17132 5160
rect 17184 5108 17190 5160
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5148 18935 5151
rect 19702 5148 19708 5160
rect 18923 5120 19708 5148
rect 18923 5117 18935 5120
rect 18877 5111 18935 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 19996 5157 20024 5188
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21192 5188 21373 5216
rect 21192 5157 21220 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5216 22431 5219
rect 22419 5188 22600 5216
rect 22419 5185 22431 5188
rect 22373 5179 22431 5185
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 20349 5151 20407 5157
rect 20349 5117 20361 5151
rect 20395 5148 20407 5151
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 20395 5120 20545 5148
rect 20395 5117 20407 5120
rect 20349 5111 20407 5117
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5148 20683 5151
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20671 5120 20821 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5148 20959 5151
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20947 5120 21097 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21085 5117 21097 5120
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 21266 5108 21272 5160
rect 21324 5108 21330 5160
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 22572 5157 22600 5188
rect 22557 5151 22615 5157
rect 22557 5117 22569 5151
rect 22603 5117 22615 5151
rect 22557 5111 22615 5117
rect 22649 5151 22707 5157
rect 22649 5117 22661 5151
rect 22695 5148 22707 5151
rect 22833 5151 22891 5157
rect 22833 5148 22845 5151
rect 22695 5120 22845 5148
rect 22695 5117 22707 5120
rect 22649 5111 22707 5117
rect 22833 5117 22845 5120
rect 22879 5117 22891 5151
rect 22833 5111 22891 5117
rect 22925 5151 22983 5157
rect 22925 5117 22937 5151
rect 22971 5148 22983 5151
rect 23109 5151 23167 5157
rect 23109 5148 23121 5151
rect 22971 5120 23121 5148
rect 22971 5117 22983 5120
rect 22925 5111 22983 5117
rect 23109 5117 23121 5120
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 23201 5151 23259 5157
rect 23201 5117 23213 5151
rect 23247 5148 23259 5151
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 23247 5120 23397 5148
rect 23247 5117 23259 5120
rect 23201 5111 23259 5117
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 23477 5151 23535 5157
rect 23477 5117 23489 5151
rect 23523 5148 23535 5151
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23523 5120 23857 5148
rect 23523 5117 23535 5120
rect 23477 5111 23535 5117
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 23845 5111 23903 5117
rect 23937 5151 23995 5157
rect 23937 5117 23949 5151
rect 23983 5148 23995 5151
rect 24121 5151 24179 5157
rect 24121 5148 24133 5151
rect 23983 5120 24133 5148
rect 23983 5117 23995 5120
rect 23937 5111 23995 5117
rect 24121 5117 24133 5120
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5148 24271 5151
rect 24397 5151 24455 5157
rect 24397 5148 24409 5151
rect 24259 5120 24409 5148
rect 24259 5117 24271 5120
rect 24213 5111 24271 5117
rect 24397 5117 24409 5120
rect 24443 5117 24455 5151
rect 24397 5111 24455 5117
rect 24489 5151 24547 5157
rect 24489 5117 24501 5151
rect 24535 5148 24547 5151
rect 24673 5151 24731 5157
rect 24673 5148 24685 5151
rect 24535 5120 24685 5148
rect 24535 5117 24547 5120
rect 24489 5111 24547 5117
rect 24673 5117 24685 5120
rect 24719 5117 24731 5151
rect 24673 5111 24731 5117
rect 24765 5151 24823 5157
rect 24765 5117 24777 5151
rect 24811 5148 24823 5151
rect 24949 5151 25007 5157
rect 24949 5148 24961 5151
rect 24811 5120 24961 5148
rect 24811 5117 24823 5120
rect 24765 5111 24823 5117
rect 24949 5117 24961 5120
rect 24995 5117 25007 5151
rect 24949 5111 25007 5117
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5117 25283 5151
rect 25225 5111 25283 5117
rect 25317 5151 25375 5157
rect 25317 5117 25329 5151
rect 25363 5148 25375 5151
rect 25501 5151 25559 5157
rect 25501 5148 25513 5151
rect 25363 5120 25513 5148
rect 25363 5117 25375 5120
rect 25317 5111 25375 5117
rect 25501 5117 25513 5120
rect 25547 5117 25559 5151
rect 25501 5111 25559 5117
rect 15197 5083 15255 5089
rect 15197 5080 15209 5083
rect 14936 5052 15209 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 15197 5049 15209 5052
rect 15243 5049 15255 5083
rect 15197 5043 15255 5049
rect 24578 5040 24584 5092
rect 24636 5080 24642 5092
rect 25240 5080 25268 5111
rect 24636 5052 25268 5080
rect 24636 5040 24642 5052
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7064 4984 7389 5012
rect 7064 4972 7070 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 7377 4975 7435 4981
rect 14918 4972 14924 5024
rect 14976 4972 14982 5024
rect 24486 4972 24492 5024
rect 24544 5012 24550 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 24544 4984 25053 5012
rect 24544 4972 24550 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 25041 4975 25099 4981
rect 25590 4972 25596 5024
rect 25648 4972 25654 5024
rect 552 4922 31648 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31648 4922
rect 552 4848 31648 4870
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 9490 4808 9496 4820
rect 8987 4780 9496 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21266 4808 21272 4820
rect 21039 4780 21272 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 24397 4811 24455 4817
rect 24397 4777 24409 4811
rect 24443 4808 24455 4811
rect 24578 4808 24584 4820
rect 24443 4780 24584 4808
rect 24443 4777 24455 4780
rect 24397 4771 24455 4777
rect 24578 4768 24584 4780
rect 24636 4768 24642 4820
rect 24946 4768 24952 4820
rect 25004 4768 25010 4820
rect 8665 4743 8723 4749
rect 8665 4709 8677 4743
rect 8711 4740 8723 4743
rect 13449 4743 13507 4749
rect 8711 4712 9444 4740
rect 8711 4709 8723 4712
rect 8665 4703 8723 4709
rect 7006 4632 7012 4684
rect 7064 4632 7070 4684
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 7239 4644 7389 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7515 4644 7665 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7116 4604 7144 4635
rect 8570 4632 8576 4684
rect 8628 4632 8634 4684
rect 9416 4681 9444 4712
rect 13449 4709 13461 4743
rect 13495 4740 13507 4743
rect 15289 4743 15347 4749
rect 13495 4712 13952 4740
rect 13495 4709 13507 4712
rect 13449 4703 13507 4709
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4672 9091 4675
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 9079 4644 9229 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 11471 4644 11621 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11882 4672 11888 4684
rect 11747 4644 11888 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 6963 4576 7144 4604
rect 9324 4604 9352 4635
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 12023 4644 12173 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 12299 4644 12449 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4672 12587 4675
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12575 4644 12725 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 12713 4641 12725 4644
rect 12759 4641 12771 4675
rect 12713 4635 12771 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12851 4644 13001 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 12989 4641 13001 4644
rect 13035 4641 13047 4675
rect 12989 4635 13047 4641
rect 13081 4675 13139 4681
rect 13081 4641 13093 4675
rect 13127 4641 13139 4675
rect 13081 4635 13139 4641
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13587 4644 13737 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9324 4576 9505 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 13096 4604 13124 4635
rect 13814 4632 13820 4684
rect 13872 4632 13878 4684
rect 13924 4681 13952 4712
rect 15289 4709 15301 4743
rect 15335 4740 15347 4743
rect 15335 4712 16160 4740
rect 15335 4709 15347 4712
rect 15289 4703 15347 4709
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4641 13967 4675
rect 13909 4635 13967 4641
rect 14918 4632 14924 4684
rect 14976 4632 14982 4684
rect 16132 4681 16160 4712
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4672 15071 4675
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 15059 4644 15209 4672
rect 15059 4641 15071 4644
rect 15013 4635 15071 4641
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 15749 4675 15807 4681
rect 15749 4641 15761 4675
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 13096 4576 14013 4604
rect 9493 4567 9551 4573
rect 14001 4573 14013 4576
rect 14047 4573 14059 4607
rect 15764 4604 15792 4635
rect 17402 4632 17408 4684
rect 17460 4632 17466 4684
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4672 17555 4675
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 17543 4644 17693 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17819 4644 17969 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 18095 4644 18245 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18233 4641 18245 4644
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 18371 4644 18521 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 18509 4641 18521 4644
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4672 18659 4675
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 18647 4644 18797 4672
rect 18647 4641 18659 4644
rect 18601 4635 18659 4641
rect 18785 4641 18797 4644
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18923 4644 19073 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4672 19211 4675
rect 19337 4675 19395 4681
rect 19337 4672 19349 4675
rect 19199 4644 19349 4672
rect 19199 4641 19211 4644
rect 19153 4635 19211 4641
rect 19337 4641 19349 4644
rect 19383 4641 19395 4675
rect 19337 4635 19395 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19475 4644 19625 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19889 4675 19947 4681
rect 19889 4672 19901 4675
rect 19751 4644 19901 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19889 4641 19901 4644
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 21085 4675 21143 4681
rect 21085 4641 21097 4675
rect 21131 4672 21143 4675
rect 21361 4675 21419 4681
rect 21361 4672 21373 4675
rect 21131 4644 21373 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 21361 4641 21373 4644
rect 21407 4641 21419 4675
rect 21361 4635 21419 4641
rect 21453 4675 21511 4681
rect 21453 4641 21465 4675
rect 21499 4672 21511 4675
rect 21637 4675 21695 4681
rect 21637 4672 21649 4675
rect 21499 4644 21649 4672
rect 21499 4641 21511 4644
rect 21453 4635 21511 4641
rect 21637 4641 21649 4644
rect 21683 4641 21695 4675
rect 21637 4635 21695 4641
rect 21729 4675 21787 4681
rect 21729 4641 21741 4675
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 16209 4607 16267 4613
rect 16209 4604 16221 4607
rect 15764 4576 16221 4604
rect 14001 4567 14059 4573
rect 16209 4573 16221 4576
rect 16255 4573 16267 4607
rect 21744 4604 21772 4635
rect 21818 4632 21824 4684
rect 21876 4632 21882 4684
rect 24486 4632 24492 4684
rect 24544 4632 24550 4684
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4672 25099 4675
rect 25590 4672 25596 4684
rect 25087 4644 25596 4672
rect 25087 4641 25099 4644
rect 25041 4635 25099 4641
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 21744 4576 21925 4604
rect 16209 4567 16267 4573
rect 21913 4573 21925 4576
rect 21959 4573 21971 4607
rect 21913 4567 21971 4573
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7745 4471 7803 4477
rect 7745 4468 7757 4471
rect 7064 4440 7757 4468
rect 7064 4428 7070 4440
rect 7745 4437 7757 4440
rect 7791 4437 7803 4471
rect 7745 4431 7803 4437
rect 11330 4428 11336 4480
rect 11388 4428 11394 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 12066 4468 12072 4480
rect 11931 4440 12072 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 15654 4428 15660 4480
rect 15712 4428 15718 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 19981 4471 20039 4477
rect 19981 4468 19993 4471
rect 19668 4440 19993 4468
rect 19668 4428 19674 4440
rect 19981 4437 19993 4440
rect 20027 4437 20039 4471
rect 19981 4431 20039 4437
rect 552 4378 31648 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31648 4378
rect 552 4304 31648 4326
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8628 4236 8677 4264
rect 8628 4224 8634 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 8665 4227 8723 4233
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11940 4236 12173 4264
rect 11940 4224 11946 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 17402 4224 17408 4276
rect 17460 4264 17466 4276
rect 17497 4267 17555 4273
rect 17497 4264 17509 4267
rect 17460 4236 17509 4264
rect 17460 4224 17466 4236
rect 17497 4233 17509 4236
rect 17543 4233 17555 4267
rect 17497 4227 17555 4233
rect 21361 4267 21419 4273
rect 21361 4233 21373 4267
rect 21407 4264 21419 4267
rect 21818 4264 21824 4276
rect 21407 4236 21824 4264
rect 21407 4233 21419 4236
rect 21361 4227 21419 4233
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 6886 4100 7481 4128
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4060 6791 4063
rect 6886 4060 6914 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8159 4100 9168 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 6779 4032 6914 4060
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 7006 4020 7012 4072
rect 7064 4020 7070 4072
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4060 7251 4063
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7239 4032 7389 4060
rect 7239 4029 7251 4032
rect 7193 4023 7251 4029
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8294 4060 8300 4072
rect 8251 4032 8300 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 6917 3995 6975 4001
rect 6917 3961 6929 3995
rect 6963 3992 6975 3995
rect 7116 3992 7144 4023
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 9140 4069 9168 4100
rect 24394 4088 24400 4140
rect 24452 4128 24458 4140
rect 24452 4100 24992 4128
rect 24452 4088 24458 4100
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4060 8815 4063
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8803 4032 8953 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10275 4032 10425 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10551 4032 10701 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10827 4032 10977 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 11103 4032 11253 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 11333 4023 11391 4029
rect 6963 3964 7144 3992
rect 9048 3992 9076 4023
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 9048 3964 9229 3992
rect 6963 3961 6975 3964
rect 6917 3955 6975 3961
rect 9217 3961 9229 3964
rect 9263 3961 9275 3995
rect 11348 3992 11376 4023
rect 11422 4020 11428 4072
rect 11480 4020 11486 4072
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4060 13967 4063
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13955 4032 14105 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14231 4032 14381 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14507 4032 14657 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14783 4032 14933 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 15059 4032 15209 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4060 15347 4063
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15335 4032 15485 4060
rect 15335 4029 15347 4032
rect 15289 4023 15347 4029
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4029 15623 4063
rect 15565 4023 15623 4029
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 11348 3964 11529 3992
rect 9217 3955 9275 3961
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 15580 3992 15608 4023
rect 15654 4020 15660 4072
rect 15712 4020 15718 4072
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4060 15807 4063
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15795 4032 15945 4060
rect 15795 4029 15807 4032
rect 15749 4023 15807 4029
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 16071 4032 16221 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4060 17647 4063
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 17635 4032 17785 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15580 3964 16313 3992
rect 11517 3955 11575 3961
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 17880 3992 17908 4023
rect 17954 4020 17960 4072
rect 18012 4020 18018 4072
rect 19610 4020 19616 4072
rect 19668 4020 19674 4072
rect 24964 4069 24992 4100
rect 19705 4063 19763 4069
rect 19705 4029 19717 4063
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19843 4032 19993 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4060 20131 4063
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 20119 4032 20269 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 21453 4063 21511 4069
rect 21453 4029 21465 4063
rect 21499 4060 21511 4063
rect 21637 4063 21695 4069
rect 21637 4060 21649 4063
rect 21499 4032 21649 4060
rect 21499 4029 21511 4032
rect 21453 4023 21511 4029
rect 21637 4029 21649 4032
rect 21683 4029 21695 4063
rect 21637 4023 21695 4029
rect 21729 4063 21787 4069
rect 21729 4029 21741 4063
rect 21775 4060 21787 4063
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 21775 4032 21925 4060
rect 21775 4029 21787 4032
rect 21729 4023 21787 4029
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22189 4063 22247 4069
rect 22189 4060 22201 4063
rect 22051 4032 22201 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22189 4029 22201 4032
rect 22235 4029 22247 4063
rect 22189 4023 22247 4029
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4060 22339 4063
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22327 4032 22477 4060
rect 22327 4029 22339 4032
rect 22281 4023 22339 4029
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 22557 4063 22615 4069
rect 22557 4029 22569 4063
rect 22603 4060 22615 4063
rect 22741 4063 22799 4069
rect 22741 4060 22753 4063
rect 22603 4032 22753 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 22741 4029 22753 4032
rect 22787 4029 22799 4063
rect 22741 4023 22799 4029
rect 22833 4063 22891 4069
rect 22833 4029 22845 4063
rect 22879 4060 22891 4063
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22879 4032 23029 4060
rect 22879 4029 22891 4032
rect 22833 4023 22891 4029
rect 23017 4029 23029 4032
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 23109 4063 23167 4069
rect 23109 4029 23121 4063
rect 23155 4060 23167 4063
rect 23293 4063 23351 4069
rect 23293 4060 23305 4063
rect 23155 4032 23305 4060
rect 23155 4029 23167 4032
rect 23109 4023 23167 4029
rect 23293 4029 23305 4032
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 23385 4063 23443 4069
rect 23385 4029 23397 4063
rect 23431 4060 23443 4063
rect 23569 4063 23627 4069
rect 23569 4060 23581 4063
rect 23431 4032 23581 4060
rect 23431 4029 23443 4032
rect 23385 4023 23443 4029
rect 23569 4029 23581 4032
rect 23615 4029 23627 4063
rect 23569 4023 23627 4029
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4060 23719 4063
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 23707 4032 23949 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 23937 4029 23949 4032
rect 23983 4029 23995 4063
rect 23937 4023 23995 4029
rect 24029 4063 24087 4069
rect 24029 4029 24041 4063
rect 24075 4060 24087 4063
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 24075 4032 24225 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4060 24363 4063
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24351 4032 24501 4060
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4060 24639 4063
rect 24765 4063 24823 4069
rect 24765 4060 24777 4063
rect 24627 4032 24777 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 24765 4029 24777 4032
rect 24811 4029 24823 4063
rect 24765 4023 24823 4029
rect 24857 4063 24915 4069
rect 24857 4029 24869 4063
rect 24903 4029 24915 4063
rect 24857 4023 24915 4029
rect 24949 4063 25007 4069
rect 24949 4029 24961 4063
rect 24995 4029 25007 4063
rect 24949 4023 25007 4029
rect 18049 3995 18107 4001
rect 18049 3992 18061 3995
rect 17880 3964 18061 3992
rect 16301 3955 16359 3961
rect 18049 3961 18061 3964
rect 18095 3961 18107 3995
rect 18049 3955 18107 3961
rect 19521 3995 19579 4001
rect 19521 3961 19533 3995
rect 19567 3992 19579 3995
rect 19720 3992 19748 4023
rect 19567 3964 19748 3992
rect 24872 3992 24900 4023
rect 25130 4020 25136 4072
rect 25188 4060 25194 4072
rect 25225 4063 25283 4069
rect 25225 4060 25237 4063
rect 25188 4032 25237 4060
rect 25188 4020 25194 4032
rect 25225 4029 25237 4032
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 25041 3995 25099 4001
rect 25041 3992 25053 3995
rect 24872 3964 25053 3992
rect 19567 3961 19579 3964
rect 19521 3955 19579 3961
rect 25041 3961 25053 3964
rect 25087 3961 25099 3995
rect 25700 3992 25728 4023
rect 25774 4020 25780 4072
rect 25832 4020 25838 4072
rect 26237 4063 26295 4069
rect 26237 4029 26249 4063
rect 26283 4060 26295 4063
rect 26421 4063 26479 4069
rect 26421 4060 26433 4063
rect 26283 4032 26433 4060
rect 26283 4029 26295 4032
rect 26237 4023 26295 4029
rect 26421 4029 26433 4032
rect 26467 4029 26479 4063
rect 26421 4023 26479 4029
rect 26513 4063 26571 4069
rect 26513 4029 26525 4063
rect 26559 4060 26571 4063
rect 26697 4063 26755 4069
rect 26697 4060 26709 4063
rect 26559 4032 26709 4060
rect 26559 4029 26571 4032
rect 26513 4023 26571 4029
rect 26697 4029 26709 4032
rect 26743 4029 26755 4063
rect 26697 4023 26755 4029
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4029 26847 4063
rect 26789 4023 26847 4029
rect 25869 3995 25927 4001
rect 25869 3992 25881 3995
rect 25700 3964 25881 3992
rect 25041 3955 25099 3961
rect 25869 3961 25881 3964
rect 25915 3961 25927 3995
rect 26804 3992 26832 4023
rect 26878 4020 26884 4072
rect 26936 4020 26942 4072
rect 26973 3995 27031 4001
rect 26973 3992 26985 3995
rect 26804 3964 26985 3992
rect 25869 3955 25927 3961
rect 26973 3961 26985 3964
rect 27019 3961 27031 3995
rect 26973 3955 27031 3961
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 10226 3924 10232 3936
rect 10183 3896 10232 3924
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 13814 3884 13820 3936
rect 13872 3884 13878 3936
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20349 3927 20407 3933
rect 20349 3924 20361 3927
rect 20312 3896 20361 3924
rect 20312 3884 20318 3896
rect 20349 3893 20361 3896
rect 20395 3893 20407 3927
rect 20349 3887 20407 3893
rect 24486 3884 24492 3936
rect 24544 3924 24550 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 24544 3896 25329 3924
rect 24544 3884 24550 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 25590 3884 25596 3936
rect 25648 3884 25654 3936
rect 26142 3884 26148 3936
rect 26200 3884 26206 3936
rect 552 3834 31648 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31648 3834
rect 552 3760 31648 3782
rect 8294 3680 8300 3732
rect 8352 3680 8358 3732
rect 13906 3680 13912 3732
rect 13964 3680 13970 3732
rect 17313 3723 17371 3729
rect 17313 3689 17325 3723
rect 17359 3720 17371 3723
rect 17954 3720 17960 3732
rect 17359 3692 17960 3720
rect 17359 3689 17371 3692
rect 17313 3683 17371 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 20441 3723 20499 3729
rect 20441 3720 20453 3723
rect 19720 3692 20453 3720
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10060 3624 10609 3652
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6871 3556 7021 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 7147 3556 7297 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3584 7435 3587
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7423 3556 7573 3584
rect 7423 3553 7435 3556
rect 7377 3547 7435 3553
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 8386 3544 8392 3596
rect 8444 3544 8450 3596
rect 10060 3593 10088 3624
rect 10597 3621 10609 3624
rect 10643 3621 10655 3655
rect 10597 3615 10655 3621
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8711 3556 8861 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8987 3556 9137 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3584 9275 3587
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 9263 3556 9413 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9401 3553 9413 3556
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9539 3556 9689 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9815 3556 9965 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10226 3544 10232 3596
rect 10284 3544 10290 3596
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 10367 3556 10517 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12676 3556 12725 3584
rect 12676 3544 12682 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 13044 3556 13277 3584
rect 13044 3544 13050 3556
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13814 3544 13820 3596
rect 13872 3544 13878 3596
rect 17405 3587 17463 3593
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17451 3556 17601 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 17589 3547 17647 3553
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3584 17739 3587
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17727 3556 17877 3584
rect 17727 3553 17739 3556
rect 17681 3547 17739 3553
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 17972 3516 18000 3547
rect 18046 3544 18052 3596
rect 18104 3544 18110 3596
rect 19720 3593 19748 3692
rect 20441 3689 20453 3692
rect 20487 3689 20499 3723
rect 20441 3683 20499 3689
rect 24394 3680 24400 3732
rect 24452 3680 24458 3732
rect 24673 3723 24731 3729
rect 24673 3689 24685 3723
rect 24719 3720 24731 3723
rect 25130 3720 25136 3732
rect 24719 3692 25136 3720
rect 24719 3689 24731 3692
rect 24673 3683 24731 3689
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 25225 3723 25283 3729
rect 25225 3689 25237 3723
rect 25271 3720 25283 3723
rect 25774 3720 25780 3732
rect 25271 3692 25780 3720
rect 25271 3689 25283 3692
rect 25225 3683 25283 3689
rect 25774 3680 25780 3692
rect 25832 3680 25838 3732
rect 26513 3723 26571 3729
rect 26513 3689 26525 3723
rect 26559 3720 26571 3723
rect 26878 3720 26884 3732
rect 26559 3692 26884 3720
rect 26559 3689 26571 3692
rect 26513 3683 26571 3689
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 20254 3652 20260 3664
rect 19996 3624 20260 3652
rect 19996 3593 20024 3624
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 25590 3652 25596 3664
rect 24780 3624 25596 3652
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3584 19487 3587
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 19475 3556 19625 3584
rect 19475 3553 19487 3556
rect 19429 3547 19487 3553
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 20073 3587 20131 3593
rect 20073 3553 20085 3587
rect 20119 3553 20131 3587
rect 20073 3547 20131 3553
rect 20165 3587 20223 3593
rect 20165 3553 20177 3587
rect 20211 3584 20223 3587
rect 20349 3587 20407 3593
rect 20349 3584 20361 3587
rect 20211 3556 20361 3584
rect 20211 3553 20223 3556
rect 20165 3547 20223 3553
rect 20349 3553 20361 3556
rect 20395 3553 20407 3587
rect 20349 3547 20407 3553
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17972 3488 18153 3516
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 20088 3516 20116 3547
rect 24486 3544 24492 3596
rect 24544 3544 24550 3596
rect 24780 3593 24808 3624
rect 25590 3612 25596 3624
rect 25648 3612 25654 3664
rect 27617 3655 27675 3661
rect 27617 3652 27629 3655
rect 27448 3624 27629 3652
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25317 3587 25375 3593
rect 25317 3553 25329 3587
rect 25363 3584 25375 3587
rect 26142 3584 26148 3596
rect 25363 3556 26148 3584
rect 25363 3553 25375 3556
rect 25317 3547 25375 3553
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 27448 3593 27476 3624
rect 27617 3621 27629 3624
rect 27663 3621 27675 3655
rect 27617 3615 27675 3621
rect 26605 3587 26663 3593
rect 26605 3553 26617 3587
rect 26651 3584 26663 3587
rect 26789 3587 26847 3593
rect 26789 3584 26801 3587
rect 26651 3556 26801 3584
rect 26651 3553 26663 3556
rect 26605 3547 26663 3553
rect 26789 3553 26801 3556
rect 26835 3553 26847 3587
rect 26789 3547 26847 3553
rect 26881 3587 26939 3593
rect 26881 3553 26893 3587
rect 26927 3584 26939 3587
rect 27065 3587 27123 3593
rect 27065 3584 27077 3587
rect 26927 3556 27077 3584
rect 26927 3553 26939 3556
rect 26881 3547 26939 3553
rect 27065 3553 27077 3556
rect 27111 3553 27123 3587
rect 27065 3547 27123 3553
rect 27157 3587 27215 3593
rect 27157 3553 27169 3587
rect 27203 3584 27215 3587
rect 27341 3587 27399 3593
rect 27341 3584 27353 3587
rect 27203 3556 27353 3584
rect 27203 3553 27215 3556
rect 27157 3547 27215 3553
rect 27341 3553 27353 3556
rect 27387 3553 27399 3587
rect 27341 3547 27399 3553
rect 27433 3587 27491 3593
rect 27433 3553 27445 3587
rect 27479 3553 27491 3587
rect 27433 3547 27491 3553
rect 27522 3544 27528 3596
rect 27580 3544 27586 3596
rect 19935 3488 20116 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7653 3383 7711 3389
rect 7653 3380 7665 3383
rect 6972 3352 7665 3380
rect 6972 3340 6978 3352
rect 7653 3349 7665 3352
rect 7699 3349 7711 3383
rect 7653 3343 7711 3349
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8662 3380 8668 3392
rect 8619 3352 8668 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 12894 3380 12900 3392
rect 12851 3352 12900 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13354 3340 13360 3392
rect 13412 3340 13418 3392
rect 19337 3383 19395 3389
rect 19337 3349 19349 3383
rect 19383 3380 19395 3383
rect 19702 3380 19708 3392
rect 19383 3352 19708 3380
rect 19383 3349 19395 3352
rect 19337 3343 19395 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 552 3290 31648 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31648 3290
rect 552 3216 31648 3238
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8444 3148 8769 3176
rect 8444 3136 8450 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 8757 3139 8815 3145
rect 12618 3136 12624 3188
rect 12676 3136 12682 3188
rect 12986 3136 12992 3188
rect 13044 3136 13050 3188
rect 17681 3179 17739 3185
rect 17681 3145 17693 3179
rect 17727 3176 17739 3179
rect 18046 3176 18052 3188
rect 17727 3148 18052 3176
rect 17727 3145 17739 3148
rect 17681 3139 17739 3145
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 26697 3179 26755 3185
rect 26697 3145 26709 3179
rect 26743 3176 26755 3179
rect 27522 3176 27528 3188
rect 26743 3148 27528 3176
rect 26743 3145 26755 3148
rect 26697 3139 26755 3145
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 19245 3111 19303 3117
rect 19245 3108 19257 3111
rect 18524 3080 19257 3108
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 7101 3043 7159 3049
rect 6595 3012 7052 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6687 2944 6837 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7024 2981 7052 3012
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 11517 3043 11575 3049
rect 7147 3012 7696 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7668 2981 7696 3012
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 15749 3043 15807 3049
rect 11563 3012 11744 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 7576 2904 7604 2935
rect 8662 2932 8668 2984
rect 8720 2932 8726 2984
rect 11054 2932 11060 2984
rect 11112 2932 11118 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 7745 2907 7803 2913
rect 7745 2904 7757 2907
rect 7576 2876 7757 2904
rect 7745 2873 7757 2876
rect 7791 2873 7803 2907
rect 7745 2867 7803 2873
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 11164 2904 11192 2935
rect 11606 2932 11612 2984
rect 11664 2932 11670 2984
rect 11716 2981 11744 3012
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 15795 3012 15976 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11839 2944 11989 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 12115 2944 12265 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2972 12403 2975
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 12391 2944 12541 2972
rect 12391 2941 12403 2944
rect 12345 2935 12403 2941
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 12894 2932 12900 2984
rect 12952 2932 12958 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13863 2944 14013 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14139 2944 14289 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14415 2944 14565 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2972 14703 2975
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14691 2944 14841 2972
rect 14691 2941 14703 2944
rect 14645 2935 14703 2941
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 11011 2876 11192 2904
rect 13740 2904 13768 2935
rect 15838 2932 15844 2984
rect 15896 2932 15902 2984
rect 15948 2981 15976 3012
rect 18524 2981 18552 3080
rect 19245 3077 19257 3080
rect 19291 3077 19303 3111
rect 19245 3071 19303 3077
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3040 19027 3043
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19015 3012 19196 3040
rect 19015 3009 19027 3012
rect 18969 3003 19027 3009
rect 19168 2981 19196 3012
rect 19628 3012 19809 3040
rect 19628 2981 19656 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3040 26479 3043
rect 26467 3012 27200 3040
rect 26467 3009 26479 3012
rect 26421 3003 26479 3009
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2941 15991 2975
rect 15933 2935 15991 2941
rect 16025 2975 16083 2981
rect 16025 2941 16037 2975
rect 16071 2972 16083 2975
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 16071 2944 16221 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 16347 2944 16497 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 16485 2941 16497 2944
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2972 16635 2975
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 16623 2944 16773 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 16761 2941 16773 2944
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16899 2944 17049 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17175 2944 17325 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 17451 2944 17601 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 17589 2935 17647 2941
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2941 19671 2975
rect 19613 2935 19671 2941
rect 19076 2904 19104 2935
rect 19702 2932 19708 2984
rect 19760 2932 19766 2984
rect 20714 2932 20720 2984
rect 20772 2932 20778 2984
rect 20809 2975 20867 2981
rect 20809 2941 20821 2975
rect 20855 2972 20867 2975
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20855 2944 21005 2972
rect 20855 2941 20867 2944
rect 20809 2935 20867 2941
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 21085 2975 21143 2981
rect 21085 2941 21097 2975
rect 21131 2972 21143 2975
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 21131 2944 21281 2972
rect 21131 2941 21143 2944
rect 21085 2935 21143 2941
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 21269 2935 21327 2941
rect 21361 2975 21419 2981
rect 21361 2941 21373 2975
rect 21407 2972 21419 2975
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 21407 2944 21557 2972
rect 21407 2941 21419 2944
rect 21361 2935 21419 2941
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21545 2935 21603 2941
rect 21637 2975 21695 2981
rect 21637 2941 21649 2975
rect 21683 2972 21695 2975
rect 21821 2975 21879 2981
rect 21821 2972 21833 2975
rect 21683 2944 21833 2972
rect 21683 2941 21695 2944
rect 21637 2935 21695 2941
rect 21821 2941 21833 2944
rect 21867 2941 21879 2975
rect 21821 2935 21879 2941
rect 21913 2975 21971 2981
rect 21913 2941 21925 2975
rect 21959 2972 21971 2975
rect 22097 2975 22155 2981
rect 22097 2972 22109 2975
rect 21959 2944 22109 2972
rect 21959 2941 21971 2944
rect 21913 2935 21971 2941
rect 22097 2941 22109 2944
rect 22143 2941 22155 2975
rect 22097 2935 22155 2941
rect 22189 2975 22247 2981
rect 22189 2941 22201 2975
rect 22235 2972 22247 2975
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 22235 2944 22385 2972
rect 22235 2941 22247 2944
rect 22189 2935 22247 2941
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22511 2944 22661 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 22741 2975 22799 2981
rect 22741 2941 22753 2975
rect 22787 2972 22799 2975
rect 22925 2975 22983 2981
rect 22925 2972 22937 2975
rect 22787 2944 22937 2972
rect 22787 2941 22799 2944
rect 22741 2935 22799 2941
rect 22925 2941 22937 2944
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 23017 2975 23075 2981
rect 23017 2941 23029 2975
rect 23063 2972 23075 2975
rect 23201 2975 23259 2981
rect 23201 2972 23213 2975
rect 23063 2944 23213 2972
rect 23063 2941 23075 2944
rect 23017 2935 23075 2941
rect 23201 2941 23213 2944
rect 23247 2941 23259 2975
rect 23201 2935 23259 2941
rect 23293 2975 23351 2981
rect 23293 2941 23305 2975
rect 23339 2972 23351 2975
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 23339 2944 23489 2972
rect 23339 2941 23351 2944
rect 23293 2935 23351 2941
rect 23477 2941 23489 2944
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 23569 2975 23627 2981
rect 23569 2941 23581 2975
rect 23615 2972 23627 2975
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23615 2944 23857 2972
rect 23615 2941 23627 2944
rect 23569 2935 23627 2941
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 23845 2935 23903 2941
rect 23937 2975 23995 2981
rect 23937 2941 23949 2975
rect 23983 2972 23995 2975
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23983 2944 24133 2972
rect 23983 2941 23995 2944
rect 23937 2935 23995 2941
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24213 2975 24271 2981
rect 24213 2941 24225 2975
rect 24259 2972 24271 2975
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 24259 2944 24409 2972
rect 24259 2941 24271 2944
rect 24213 2935 24271 2941
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 26510 2932 26516 2984
rect 26568 2932 26574 2984
rect 27172 2981 27200 3012
rect 26789 2975 26847 2981
rect 26789 2941 26801 2975
rect 26835 2972 26847 2975
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26835 2944 26985 2972
rect 26835 2941 26847 2944
rect 26789 2935 26847 2941
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27065 2975 27123 2981
rect 27065 2941 27077 2975
rect 27111 2941 27123 2975
rect 27065 2935 27123 2941
rect 27157 2975 27215 2981
rect 27157 2941 27169 2975
rect 27203 2941 27215 2975
rect 27157 2935 27215 2941
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 13740 2876 13860 2904
rect 19076 2876 19533 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 13832 2848 13860 2876
rect 19521 2873 19533 2876
rect 19567 2873 19579 2907
rect 27080 2904 27108 2935
rect 27249 2907 27307 2913
rect 27249 2904 27261 2907
rect 27080 2876 27261 2904
rect 19521 2867 19579 2873
rect 27249 2873 27261 2876
rect 27295 2873 27307 2907
rect 27249 2867 27307 2873
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7558 2836 7564 2848
rect 7515 2808 7564 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 11698 2836 11704 2848
rect 11287 2808 11704 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 13265 2839 13323 2845
rect 13265 2805 13277 2839
rect 13311 2836 13323 2839
rect 13722 2836 13728 2848
rect 13311 2808 13728 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 13814 2796 13820 2848
rect 13872 2796 13878 2848
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 14332 2808 14933 2836
rect 14332 2796 14338 2808
rect 14921 2805 14933 2808
rect 14967 2805 14979 2839
rect 14921 2799 14979 2805
rect 18417 2839 18475 2845
rect 18417 2805 18429 2839
rect 18463 2836 18475 2839
rect 18782 2836 18788 2848
rect 18463 2808 18788 2836
rect 18463 2805 18475 2808
rect 18417 2799 18475 2805
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 23934 2796 23940 2848
rect 23992 2836 23998 2848
rect 24489 2839 24547 2845
rect 24489 2836 24501 2839
rect 23992 2808 24501 2836
rect 23992 2796 23998 2808
rect 24489 2805 24501 2808
rect 24535 2805 24547 2839
rect 24489 2799 24547 2805
rect 552 2746 31648 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31648 2746
rect 552 2672 31648 2694
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 11112 2604 11253 2632
rect 11112 2592 11118 2604
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 11241 2595 11299 2601
rect 11606 2592 11612 2644
rect 11664 2632 11670 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 11664 2604 11805 2632
rect 11664 2592 11670 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 11793 2595 11851 2601
rect 13814 2592 13820 2644
rect 13872 2592 13878 2644
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 9401 2567 9459 2573
rect 9401 2564 9413 2567
rect 8956 2536 9413 2564
rect 7558 2456 7564 2508
rect 7616 2456 7622 2508
rect 8956 2505 8984 2536
rect 9401 2533 9413 2536
rect 9447 2533 9459 2567
rect 9401 2527 9459 2533
rect 10689 2567 10747 2573
rect 10689 2533 10701 2567
rect 10735 2564 10747 2567
rect 14185 2567 14243 2573
rect 10735 2536 11468 2564
rect 10735 2533 10747 2536
rect 10689 2527 10747 2533
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7699 2468 7849 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2496 7987 2499
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 7975 2468 8125 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 8251 2468 8401 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2465 10563 2499
rect 10505 2459 10563 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 11054 2496 11060 2508
rect 10827 2468 11060 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2428 8907 2431
rect 9048 2428 9076 2459
rect 8895 2400 9076 2428
rect 8895 2397 8907 2400
rect 8849 2391 8907 2397
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 9324 2360 9352 2459
rect 10520 2428 10548 2459
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11440 2505 11468 2536
rect 14185 2533 14197 2567
rect 14231 2564 14243 2567
rect 15580 2564 15608 2595
rect 15838 2592 15844 2644
rect 15896 2592 15902 2644
rect 20714 2592 20720 2644
rect 20772 2592 20778 2644
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 27065 2635 27123 2641
rect 27065 2632 27077 2635
rect 26568 2604 27077 2632
rect 26568 2592 26574 2604
rect 27065 2601 27077 2604
rect 27111 2601 27123 2635
rect 27065 2595 27123 2601
rect 20441 2567 20499 2573
rect 14231 2536 14412 2564
rect 15580 2536 16436 2564
rect 14231 2533 14243 2536
rect 14185 2527 14243 2533
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 11238 2428 11244 2440
rect 10520 2400 11244 2428
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11348 2428 11376 2459
rect 11698 2456 11704 2508
rect 11756 2456 11762 2508
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11348 2400 11529 2428
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 13648 2428 13676 2459
rect 13722 2456 13728 2508
rect 13780 2456 13786 2508
rect 14274 2456 14280 2508
rect 14332 2456 14338 2508
rect 14384 2505 14412 2536
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2465 14427 2499
rect 14369 2459 14427 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15562 2496 15568 2508
rect 15519 2468 15568 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 16408 2505 16436 2536
rect 20441 2533 20453 2567
rect 20487 2564 20499 2567
rect 23845 2567 23903 2573
rect 20487 2536 21312 2564
rect 20487 2533 20499 2536
rect 20441 2527 20499 2533
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 15979 2468 16221 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 16393 2499 16451 2505
rect 16393 2465 16405 2499
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13648 2400 14473 2428
rect 11517 2391 11575 2397
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 16316 2428 16344 2459
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16316 2400 16497 2428
rect 14461 2391 14519 2397
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 18708 2428 18736 2459
rect 18782 2456 18788 2508
rect 18840 2456 18846 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18923 2468 19073 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19153 2499 19211 2505
rect 19153 2465 19165 2499
rect 19199 2496 19211 2499
rect 19337 2499 19395 2505
rect 19337 2496 19349 2499
rect 19199 2468 19349 2496
rect 19199 2465 19211 2468
rect 19153 2459 19211 2465
rect 19337 2465 19349 2468
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 20533 2499 20591 2505
rect 20533 2465 20545 2499
rect 20579 2496 20591 2499
rect 20622 2496 20628 2508
rect 20579 2468 20628 2496
rect 20579 2465 20591 2468
rect 20533 2459 20591 2465
rect 20622 2456 20628 2468
rect 20680 2456 20686 2508
rect 21284 2505 21312 2536
rect 23845 2533 23857 2567
rect 23891 2564 23903 2567
rect 23891 2536 24072 2564
rect 23891 2533 23903 2536
rect 23845 2527 23903 2533
rect 20809 2499 20867 2505
rect 20809 2465 20821 2499
rect 20855 2496 20867 2499
rect 20993 2499 21051 2505
rect 20993 2496 21005 2499
rect 20855 2468 21005 2496
rect 20855 2465 20867 2468
rect 20809 2459 20867 2465
rect 20993 2465 21005 2468
rect 21039 2465 21051 2499
rect 20993 2459 21051 2465
rect 21085 2499 21143 2505
rect 21085 2465 21097 2499
rect 21131 2465 21143 2499
rect 21085 2459 21143 2465
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18708 2400 19441 2428
rect 16485 2391 16543 2397
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 21100 2428 21128 2459
rect 23934 2456 23940 2508
rect 23992 2456 23998 2508
rect 24044 2505 24072 2536
rect 24029 2499 24087 2505
rect 24029 2465 24041 2499
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2496 24179 2499
rect 24305 2499 24363 2505
rect 24305 2496 24317 2499
rect 24167 2468 24317 2496
rect 24167 2465 24179 2468
rect 24121 2459 24179 2465
rect 24305 2465 24317 2468
rect 24351 2465 24363 2499
rect 24305 2459 24363 2465
rect 24397 2499 24455 2505
rect 24397 2465 24409 2499
rect 24443 2496 24455 2499
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24443 2468 24593 2496
rect 24443 2465 24455 2468
rect 24397 2459 24455 2465
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 24673 2499 24731 2505
rect 24673 2465 24685 2499
rect 24719 2496 24731 2499
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24719 2468 24869 2496
rect 24719 2465 24731 2468
rect 24673 2459 24731 2465
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 24949 2499 25007 2505
rect 24949 2465 24961 2499
rect 24995 2496 25007 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24995 2468 25145 2496
rect 24995 2465 25007 2468
rect 24949 2459 25007 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 25225 2499 25283 2505
rect 25225 2465 25237 2499
rect 25271 2496 25283 2499
rect 25409 2499 25467 2505
rect 25409 2496 25421 2499
rect 25271 2468 25421 2496
rect 25271 2465 25283 2468
rect 25225 2459 25283 2465
rect 25409 2465 25421 2468
rect 25455 2465 25467 2499
rect 25409 2459 25467 2465
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2496 25559 2499
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25547 2468 25697 2496
rect 25547 2465 25559 2468
rect 25501 2459 25559 2465
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 25777 2499 25835 2505
rect 25777 2465 25789 2499
rect 25823 2496 25835 2499
rect 25961 2499 26019 2505
rect 25961 2496 25973 2499
rect 25823 2468 25973 2496
rect 25823 2465 25835 2468
rect 25777 2459 25835 2465
rect 25961 2465 25973 2468
rect 26007 2465 26019 2499
rect 25961 2459 26019 2465
rect 26053 2499 26111 2505
rect 26053 2465 26065 2499
rect 26099 2496 26111 2499
rect 26421 2499 26479 2505
rect 26421 2496 26433 2499
rect 26099 2468 26433 2496
rect 26099 2465 26111 2468
rect 26053 2459 26111 2465
rect 26421 2465 26433 2468
rect 26467 2465 26479 2499
rect 26421 2459 26479 2465
rect 26513 2499 26571 2505
rect 26513 2465 26525 2499
rect 26559 2496 26571 2499
rect 26697 2499 26755 2505
rect 26697 2496 26709 2499
rect 26559 2468 26709 2496
rect 26559 2465 26571 2468
rect 26513 2459 26571 2465
rect 26697 2465 26709 2468
rect 26743 2465 26755 2499
rect 26697 2459 26755 2465
rect 26789 2499 26847 2505
rect 26789 2465 26801 2499
rect 26835 2496 26847 2499
rect 26973 2499 27031 2505
rect 26973 2496 26985 2499
rect 26835 2468 26985 2496
rect 26835 2465 26847 2468
rect 26789 2459 26847 2465
rect 26973 2465 26985 2468
rect 27019 2465 27031 2499
rect 26973 2459 27031 2465
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21100 2400 21373 2428
rect 19429 2391 19487 2397
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 8527 2332 9352 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 9088 2264 9137 2292
rect 9088 2252 9094 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 10410 2252 10416 2304
rect 10468 2252 10474 2304
rect 13538 2252 13544 2304
rect 13596 2252 13602 2304
rect 18598 2252 18604 2304
rect 18656 2252 18662 2304
rect 552 2202 31648 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31648 2202
rect 552 2128 31648 2150
rect 11054 2048 11060 2100
rect 11112 2048 11118 2100
rect 11238 2048 11244 2100
rect 11296 2088 11302 2100
rect 11333 2091 11391 2097
rect 11333 2088 11345 2091
rect 11296 2060 11345 2088
rect 11296 2048 11302 2060
rect 11333 2057 11345 2060
rect 11379 2057 11391 2091
rect 11333 2051 11391 2057
rect 15562 2048 15568 2100
rect 15620 2048 15626 2100
rect 20622 2048 20628 2100
rect 20680 2048 20686 2100
rect 10781 2023 10839 2029
rect 10781 1989 10793 2023
rect 10827 2020 10839 2023
rect 10827 1992 11836 2020
rect 10827 1989 10839 1992
rect 10781 1983 10839 1989
rect 8941 1955 8999 1961
rect 8941 1921 8953 1955
rect 8987 1952 8999 1955
rect 8987 1924 9168 1952
rect 8987 1921 8999 1924
rect 8941 1915 8999 1921
rect 8757 1887 8815 1893
rect 8757 1853 8769 1887
rect 8803 1853 8815 1887
rect 8757 1847 8815 1853
rect 8772 1816 8800 1847
rect 9030 1844 9036 1896
rect 9088 1844 9094 1896
rect 9140 1893 9168 1924
rect 10410 1912 10416 1964
rect 10468 1952 10474 1964
rect 10468 1924 11008 1952
rect 10468 1912 10474 1924
rect 9125 1887 9183 1893
rect 9125 1853 9137 1887
rect 9171 1853 9183 1887
rect 9125 1847 9183 1853
rect 9217 1887 9275 1893
rect 9217 1853 9229 1887
rect 9263 1884 9275 1887
rect 9401 1887 9459 1893
rect 9401 1884 9413 1887
rect 9263 1856 9413 1884
rect 9263 1853 9275 1856
rect 9217 1847 9275 1853
rect 9401 1853 9413 1856
rect 9447 1853 9459 1887
rect 9401 1847 9459 1853
rect 10870 1844 10876 1896
rect 10928 1844 10934 1896
rect 10980 1893 11008 1924
rect 11808 1893 11836 1992
rect 13909 1955 13967 1961
rect 13909 1952 13921 1955
rect 13372 1924 13921 1952
rect 13372 1893 13400 1924
rect 13909 1921 13921 1924
rect 13955 1921 13967 1955
rect 16393 1955 16451 1961
rect 16393 1952 16405 1955
rect 13909 1915 13967 1921
rect 16224 1924 16405 1952
rect 10965 1887 11023 1893
rect 10965 1853 10977 1887
rect 11011 1853 11023 1887
rect 10965 1847 11023 1853
rect 11425 1887 11483 1893
rect 11425 1853 11437 1887
rect 11471 1884 11483 1887
rect 11609 1887 11667 1893
rect 11609 1884 11621 1887
rect 11471 1856 11621 1884
rect 11471 1853 11483 1856
rect 11425 1847 11483 1853
rect 11609 1853 11621 1856
rect 11655 1853 11667 1887
rect 11609 1847 11667 1853
rect 11701 1887 11759 1893
rect 11701 1853 11713 1887
rect 11747 1853 11759 1887
rect 11701 1847 11759 1853
rect 11793 1887 11851 1893
rect 11793 1853 11805 1887
rect 11839 1853 11851 1887
rect 11793 1847 11851 1853
rect 12805 1887 12863 1893
rect 12805 1853 12817 1887
rect 12851 1884 12863 1887
rect 12989 1887 13047 1893
rect 12989 1884 13001 1887
rect 12851 1856 13001 1884
rect 12851 1853 12863 1856
rect 12805 1847 12863 1853
rect 12989 1853 13001 1856
rect 13035 1853 13047 1887
rect 12989 1847 13047 1853
rect 13081 1887 13139 1893
rect 13081 1853 13093 1887
rect 13127 1884 13139 1887
rect 13265 1887 13323 1893
rect 13265 1884 13277 1887
rect 13127 1856 13277 1884
rect 13127 1853 13139 1856
rect 13081 1847 13139 1853
rect 13265 1853 13277 1856
rect 13311 1853 13323 1887
rect 13265 1847 13323 1853
rect 13357 1887 13415 1893
rect 13357 1853 13369 1887
rect 13403 1853 13415 1887
rect 13357 1847 13415 1853
rect 9493 1819 9551 1825
rect 9493 1816 9505 1819
rect 8772 1788 9505 1816
rect 9493 1785 9505 1788
rect 9539 1785 9551 1819
rect 11716 1816 11744 1847
rect 13538 1844 13544 1896
rect 13596 1844 13602 1896
rect 16224 1893 16252 1924
rect 16393 1921 16405 1924
rect 16439 1921 16451 1955
rect 16393 1915 16451 1921
rect 17221 1955 17279 1961
rect 17221 1921 17233 1955
rect 17267 1952 17279 1955
rect 19337 1955 19395 1961
rect 19337 1952 19349 1955
rect 17267 1924 17724 1952
rect 17267 1921 17279 1924
rect 17221 1915 17279 1921
rect 13633 1887 13691 1893
rect 13633 1853 13645 1887
rect 13679 1884 13691 1887
rect 13817 1887 13875 1893
rect 13817 1884 13829 1887
rect 13679 1856 13829 1884
rect 13679 1853 13691 1856
rect 13633 1847 13691 1853
rect 13817 1853 13829 1856
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 15657 1887 15715 1893
rect 15657 1853 15669 1887
rect 15703 1884 15715 1887
rect 15841 1887 15899 1893
rect 15841 1884 15853 1887
rect 15703 1856 15853 1884
rect 15703 1853 15715 1856
rect 15657 1847 15715 1853
rect 15841 1853 15853 1856
rect 15887 1853 15899 1887
rect 15841 1847 15899 1853
rect 15933 1887 15991 1893
rect 15933 1853 15945 1887
rect 15979 1884 15991 1887
rect 16117 1887 16175 1893
rect 16117 1884 16129 1887
rect 15979 1856 16129 1884
rect 15979 1853 15991 1856
rect 15933 1847 15991 1853
rect 16117 1853 16129 1856
rect 16163 1853 16175 1887
rect 16117 1847 16175 1853
rect 16209 1887 16267 1893
rect 16209 1853 16221 1887
rect 16255 1853 16267 1887
rect 16209 1847 16267 1853
rect 16298 1844 16304 1896
rect 16356 1844 16362 1896
rect 17696 1893 17724 1924
rect 19168 1924 19349 1952
rect 19168 1893 19196 1924
rect 19337 1921 19349 1924
rect 19383 1921 19395 1955
rect 19337 1915 19395 1921
rect 21082 1912 21088 1964
rect 21140 1952 21146 1964
rect 21140 1924 21404 1952
rect 21140 1912 21146 1924
rect 21376 1893 21404 1924
rect 17313 1887 17371 1893
rect 17313 1853 17325 1887
rect 17359 1884 17371 1887
rect 17497 1887 17555 1893
rect 17497 1884 17509 1887
rect 17359 1856 17509 1884
rect 17359 1853 17371 1856
rect 17313 1847 17371 1853
rect 17497 1853 17509 1856
rect 17543 1853 17555 1887
rect 17497 1847 17555 1853
rect 17589 1887 17647 1893
rect 17589 1853 17601 1887
rect 17635 1853 17647 1887
rect 17589 1847 17647 1853
rect 17681 1887 17739 1893
rect 17681 1853 17693 1887
rect 17727 1853 17739 1887
rect 17681 1847 17739 1853
rect 18141 1887 18199 1893
rect 18141 1853 18153 1887
rect 18187 1884 18199 1887
rect 18325 1887 18383 1893
rect 18325 1884 18337 1887
rect 18187 1856 18337 1884
rect 18187 1853 18199 1856
rect 18141 1847 18199 1853
rect 18325 1853 18337 1856
rect 18371 1853 18383 1887
rect 18325 1847 18383 1853
rect 18417 1887 18475 1893
rect 18417 1853 18429 1887
rect 18463 1884 18475 1887
rect 18785 1887 18843 1893
rect 18785 1884 18797 1887
rect 18463 1856 18797 1884
rect 18463 1853 18475 1856
rect 18417 1847 18475 1853
rect 18785 1853 18797 1856
rect 18831 1853 18843 1887
rect 18785 1847 18843 1853
rect 18877 1887 18935 1893
rect 18877 1853 18889 1887
rect 18923 1884 18935 1887
rect 19061 1887 19119 1893
rect 19061 1884 19073 1887
rect 18923 1856 19073 1884
rect 18923 1853 18935 1856
rect 18877 1847 18935 1853
rect 19061 1853 19073 1856
rect 19107 1853 19119 1887
rect 19061 1847 19119 1853
rect 19153 1887 19211 1893
rect 19153 1853 19165 1887
rect 19199 1853 19211 1887
rect 19153 1847 19211 1853
rect 19245 1887 19303 1893
rect 19245 1853 19257 1887
rect 19291 1853 19303 1887
rect 19245 1847 19303 1853
rect 20717 1887 20775 1893
rect 20717 1853 20729 1887
rect 20763 1884 20775 1887
rect 20901 1887 20959 1893
rect 20901 1884 20913 1887
rect 20763 1856 20913 1884
rect 20763 1853 20775 1856
rect 20717 1847 20775 1853
rect 20901 1853 20913 1856
rect 20947 1853 20959 1887
rect 20901 1847 20959 1853
rect 20993 1887 21051 1893
rect 20993 1853 21005 1887
rect 21039 1884 21051 1887
rect 21177 1887 21235 1893
rect 21177 1884 21189 1887
rect 21039 1856 21189 1884
rect 21039 1853 21051 1856
rect 20993 1847 21051 1853
rect 21177 1853 21189 1856
rect 21223 1853 21235 1887
rect 21177 1847 21235 1853
rect 21269 1887 21327 1893
rect 21269 1853 21281 1887
rect 21315 1853 21327 1887
rect 21269 1847 21327 1853
rect 21361 1887 21419 1893
rect 21361 1853 21373 1887
rect 21407 1853 21419 1887
rect 21361 1847 21419 1853
rect 11885 1819 11943 1825
rect 11885 1816 11897 1819
rect 11716 1788 11897 1816
rect 9493 1779 9551 1785
rect 11885 1785 11897 1788
rect 11931 1785 11943 1819
rect 17604 1816 17632 1847
rect 18049 1819 18107 1825
rect 18049 1816 18061 1819
rect 17604 1788 18061 1816
rect 11885 1779 11943 1785
rect 18049 1785 18061 1788
rect 18095 1785 18107 1819
rect 18049 1779 18107 1785
rect 18598 1776 18604 1828
rect 18656 1816 18662 1828
rect 19260 1816 19288 1847
rect 18656 1788 19288 1816
rect 21284 1816 21312 1847
rect 21453 1819 21511 1825
rect 21453 1816 21465 1819
rect 21284 1788 21465 1816
rect 18656 1776 18662 1788
rect 21453 1785 21465 1788
rect 21499 1785 21511 1819
rect 21453 1779 21511 1785
rect 8662 1708 8668 1760
rect 8720 1708 8726 1760
rect 12713 1751 12771 1757
rect 12713 1717 12725 1751
rect 12759 1748 12771 1751
rect 13170 1748 13176 1760
rect 12759 1720 13176 1748
rect 12759 1717 12771 1720
rect 12713 1711 12771 1717
rect 13170 1708 13176 1720
rect 13228 1708 13234 1760
rect 17218 1708 17224 1760
rect 17276 1748 17282 1760
rect 17773 1751 17831 1757
rect 17773 1748 17785 1751
rect 17276 1720 17785 1748
rect 17276 1708 17282 1720
rect 17773 1717 17785 1720
rect 17819 1717 17831 1751
rect 17773 1711 17831 1717
rect 552 1658 31648 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31648 1658
rect 552 1584 31648 1606
rect 10870 1504 10876 1556
rect 10928 1544 10934 1556
rect 11149 1547 11207 1553
rect 11149 1544 11161 1547
rect 10928 1516 11161 1544
rect 10928 1504 10934 1516
rect 11149 1513 11161 1516
rect 11195 1513 11207 1547
rect 11149 1507 11207 1513
rect 15657 1547 15715 1553
rect 15657 1513 15669 1547
rect 15703 1544 15715 1547
rect 16298 1544 16304 1556
rect 15703 1516 16304 1544
rect 15703 1513 15715 1516
rect 15657 1507 15715 1513
rect 16298 1504 16304 1516
rect 16356 1504 16362 1556
rect 20625 1547 20683 1553
rect 20625 1513 20637 1547
rect 20671 1544 20683 1547
rect 20671 1516 21772 1544
rect 20671 1513 20683 1516
rect 20625 1507 20683 1513
rect 9585 1479 9643 1485
rect 9585 1476 9597 1479
rect 9416 1448 9597 1476
rect 8662 1368 8668 1420
rect 8720 1368 8726 1420
rect 9416 1417 9444 1448
rect 9585 1445 9597 1448
rect 9631 1445 9643 1479
rect 9585 1439 9643 1445
rect 10137 1479 10195 1485
rect 10137 1445 10149 1479
rect 10183 1476 10195 1479
rect 11701 1479 11759 1485
rect 11701 1476 11713 1479
rect 10183 1448 10364 1476
rect 10183 1445 10195 1448
rect 10137 1439 10195 1445
rect 8757 1411 8815 1417
rect 8757 1377 8769 1411
rect 8803 1408 8815 1411
rect 8941 1411 8999 1417
rect 8941 1408 8953 1411
rect 8803 1380 8953 1408
rect 8803 1377 8815 1380
rect 8757 1371 8815 1377
rect 8941 1377 8953 1380
rect 8987 1377 8999 1411
rect 8941 1371 8999 1377
rect 9033 1411 9091 1417
rect 9033 1377 9045 1411
rect 9079 1408 9091 1411
rect 9401 1411 9459 1417
rect 9079 1380 9352 1408
rect 9079 1377 9091 1380
rect 9033 1371 9091 1377
rect 9324 1340 9352 1380
rect 9401 1377 9413 1411
rect 9447 1377 9459 1411
rect 9401 1371 9459 1377
rect 9493 1411 9551 1417
rect 9493 1377 9505 1411
rect 9539 1377 9551 1411
rect 9493 1371 9551 1377
rect 9508 1340 9536 1371
rect 10226 1368 10232 1420
rect 10284 1368 10290 1420
rect 10336 1417 10364 1448
rect 11532 1448 11713 1476
rect 11532 1417 11560 1448
rect 11701 1445 11713 1448
rect 11747 1445 11759 1479
rect 16485 1479 16543 1485
rect 16485 1476 16497 1479
rect 11701 1439 11759 1445
rect 16316 1448 16497 1476
rect 10321 1411 10379 1417
rect 10321 1377 10333 1411
rect 10367 1377 10379 1411
rect 10321 1371 10379 1377
rect 10413 1411 10471 1417
rect 10413 1377 10425 1411
rect 10459 1408 10471 1411
rect 10597 1411 10655 1417
rect 10597 1408 10609 1411
rect 10459 1380 10609 1408
rect 10459 1377 10471 1380
rect 10413 1371 10471 1377
rect 10597 1377 10609 1380
rect 10643 1377 10655 1411
rect 10597 1371 10655 1377
rect 10689 1411 10747 1417
rect 10689 1377 10701 1411
rect 10735 1408 10747 1411
rect 11241 1411 11299 1417
rect 10735 1380 11192 1408
rect 10735 1377 10747 1380
rect 10689 1371 10747 1377
rect 9324 1312 9536 1340
rect 11164 1340 11192 1380
rect 11241 1377 11253 1411
rect 11287 1408 11299 1411
rect 11425 1411 11483 1417
rect 11425 1408 11437 1411
rect 11287 1380 11437 1408
rect 11287 1377 11299 1380
rect 11241 1371 11299 1377
rect 11425 1377 11437 1380
rect 11471 1377 11483 1411
rect 11425 1371 11483 1377
rect 11517 1411 11575 1417
rect 11517 1377 11529 1411
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11609 1411 11667 1417
rect 11609 1377 11621 1411
rect 11655 1377 11667 1411
rect 11609 1371 11667 1377
rect 11624 1340 11652 1371
rect 13170 1368 13176 1420
rect 13228 1368 13234 1420
rect 16316 1417 16344 1448
rect 16485 1445 16497 1448
rect 16531 1445 16543 1479
rect 16485 1439 16543 1445
rect 17129 1479 17187 1485
rect 17129 1445 17141 1479
rect 17175 1476 17187 1479
rect 20901 1479 20959 1485
rect 17175 1448 17356 1476
rect 17175 1445 17187 1448
rect 17129 1439 17187 1445
rect 13265 1411 13323 1417
rect 13265 1377 13277 1411
rect 13311 1408 13323 1411
rect 13449 1411 13507 1417
rect 13449 1408 13461 1411
rect 13311 1380 13461 1408
rect 13311 1377 13323 1380
rect 13265 1371 13323 1377
rect 13449 1377 13461 1380
rect 13495 1377 13507 1411
rect 13449 1371 13507 1377
rect 13541 1411 13599 1417
rect 13541 1377 13553 1411
rect 13587 1408 13599 1411
rect 13725 1411 13783 1417
rect 13725 1408 13737 1411
rect 13587 1380 13737 1408
rect 13587 1377 13599 1380
rect 13541 1371 13599 1377
rect 13725 1377 13737 1380
rect 13771 1377 13783 1411
rect 13725 1371 13783 1377
rect 13817 1411 13875 1417
rect 13817 1377 13829 1411
rect 13863 1408 13875 1411
rect 14001 1411 14059 1417
rect 14001 1408 14013 1411
rect 13863 1380 14013 1408
rect 13863 1377 13875 1380
rect 13817 1371 13875 1377
rect 14001 1377 14013 1380
rect 14047 1377 14059 1411
rect 14001 1371 14059 1377
rect 15749 1411 15807 1417
rect 15749 1377 15761 1411
rect 15795 1408 15807 1411
rect 16209 1411 16267 1417
rect 16209 1408 16221 1411
rect 15795 1380 16221 1408
rect 15795 1377 15807 1380
rect 15749 1371 15807 1377
rect 16209 1377 16221 1380
rect 16255 1377 16267 1411
rect 16209 1371 16267 1377
rect 16301 1411 16359 1417
rect 16301 1377 16313 1411
rect 16347 1377 16359 1411
rect 16301 1371 16359 1377
rect 16390 1368 16396 1420
rect 16448 1368 16454 1420
rect 17218 1368 17224 1420
rect 17276 1368 17282 1420
rect 17328 1417 17356 1448
rect 20901 1445 20913 1479
rect 20947 1476 20959 1479
rect 21082 1476 21088 1488
rect 20947 1448 21088 1476
rect 20947 1445 20959 1448
rect 20901 1439 20959 1445
rect 21082 1436 21088 1448
rect 21140 1436 21146 1488
rect 21637 1479 21695 1485
rect 21637 1476 21649 1479
rect 21468 1448 21649 1476
rect 17313 1411 17371 1417
rect 17313 1377 17325 1411
rect 17359 1377 17371 1411
rect 17313 1371 17371 1377
rect 17405 1411 17463 1417
rect 17405 1377 17417 1411
rect 17451 1408 17463 1411
rect 17589 1411 17647 1417
rect 17589 1408 17601 1411
rect 17451 1380 17601 1408
rect 17451 1377 17463 1380
rect 17405 1371 17463 1377
rect 17589 1377 17601 1380
rect 17635 1377 17647 1411
rect 17589 1371 17647 1377
rect 18690 1368 18696 1420
rect 18748 1368 18754 1420
rect 18785 1411 18843 1417
rect 18785 1377 18797 1411
rect 18831 1408 18843 1411
rect 18969 1411 19027 1417
rect 18969 1408 18981 1411
rect 18831 1380 18981 1408
rect 18831 1377 18843 1380
rect 18785 1371 18843 1377
rect 18969 1377 18981 1380
rect 19015 1377 19027 1411
rect 18969 1371 19027 1377
rect 19061 1411 19119 1417
rect 19061 1377 19073 1411
rect 19107 1408 19119 1411
rect 19245 1411 19303 1417
rect 19245 1408 19257 1411
rect 19107 1380 19257 1408
rect 19107 1377 19119 1380
rect 19061 1371 19119 1377
rect 19245 1377 19257 1380
rect 19291 1377 19303 1411
rect 19245 1371 19303 1377
rect 19337 1411 19395 1417
rect 19337 1377 19349 1411
rect 19383 1408 19395 1411
rect 19521 1411 19579 1417
rect 19521 1408 19533 1411
rect 19383 1380 19533 1408
rect 19383 1377 19395 1380
rect 19337 1371 19395 1377
rect 19521 1377 19533 1380
rect 19567 1377 19579 1411
rect 19521 1371 19579 1377
rect 19613 1411 19671 1417
rect 19613 1377 19625 1411
rect 19659 1408 19671 1411
rect 19797 1411 19855 1417
rect 19797 1408 19809 1411
rect 19659 1380 19809 1408
rect 19659 1377 19671 1380
rect 19613 1371 19671 1377
rect 19797 1377 19809 1380
rect 19843 1377 19855 1411
rect 19797 1371 19855 1377
rect 20714 1368 20720 1420
rect 20772 1368 20778 1420
rect 21468 1417 21496 1448
rect 21637 1445 21649 1448
rect 21683 1445 21695 1479
rect 21637 1439 21695 1445
rect 20993 1411 21051 1417
rect 20993 1377 21005 1411
rect 21039 1408 21051 1411
rect 21361 1411 21419 1417
rect 21361 1408 21373 1411
rect 21039 1380 21373 1408
rect 21039 1377 21051 1380
rect 20993 1371 21051 1377
rect 21361 1377 21373 1380
rect 21407 1377 21419 1411
rect 21361 1371 21419 1377
rect 21453 1411 21511 1417
rect 21453 1377 21465 1411
rect 21499 1377 21511 1411
rect 21453 1371 21511 1377
rect 21545 1411 21603 1417
rect 21545 1377 21557 1411
rect 21591 1408 21603 1411
rect 21744 1408 21772 1516
rect 21591 1380 21772 1408
rect 21591 1377 21603 1380
rect 21545 1371 21603 1377
rect 11164 1312 11652 1340
rect 8938 1164 8944 1216
rect 8996 1204 9002 1216
rect 9309 1207 9367 1213
rect 9309 1204 9321 1207
rect 8996 1176 9321 1204
rect 8996 1164 9002 1176
rect 9309 1173 9321 1176
rect 9355 1173 9367 1207
rect 9309 1167 9367 1173
rect 13906 1164 13912 1216
rect 13964 1204 13970 1216
rect 14093 1207 14151 1213
rect 14093 1204 14105 1207
rect 13964 1176 14105 1204
rect 13964 1164 13970 1176
rect 14093 1173 14105 1176
rect 14139 1173 14151 1207
rect 14093 1167 14151 1173
rect 17310 1164 17316 1216
rect 17368 1204 17374 1216
rect 17681 1207 17739 1213
rect 17681 1204 17693 1207
rect 17368 1176 17693 1204
rect 17368 1164 17374 1176
rect 17681 1173 17693 1176
rect 17727 1173 17739 1207
rect 17681 1167 17739 1173
rect 19886 1164 19892 1216
rect 19944 1164 19950 1216
rect 552 1114 31648 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31648 1114
rect 552 1040 31648 1062
rect 10226 960 10232 1012
rect 10284 1000 10290 1012
rect 10413 1003 10471 1009
rect 10413 1000 10425 1003
rect 10284 972 10425 1000
rect 10284 960 10290 972
rect 10413 969 10425 972
rect 10459 969 10471 1003
rect 10413 963 10471 969
rect 15565 1003 15623 1009
rect 15565 969 15577 1003
rect 15611 1000 15623 1003
rect 16390 1000 16396 1012
rect 15611 972 16396 1000
rect 15611 969 15623 972
rect 15565 963 15623 969
rect 16390 960 16396 972
rect 16448 960 16454 1012
rect 18690 960 18696 1012
rect 18748 1000 18754 1012
rect 18785 1003 18843 1009
rect 18785 1000 18797 1003
rect 18748 972 18797 1000
rect 18748 960 18754 972
rect 18785 969 18797 972
rect 18831 969 18843 1003
rect 18785 963 18843 969
rect 20714 960 20720 1012
rect 20772 1000 20778 1012
rect 20993 1003 21051 1009
rect 20993 1000 21005 1003
rect 20772 972 21005 1000
rect 20772 960 20778 972
rect 20993 969 21005 972
rect 21039 969 21051 1003
rect 20993 963 21051 969
rect 8849 867 8907 873
rect 8849 833 8861 867
rect 8895 864 8907 867
rect 9953 867 10011 873
rect 8895 836 9076 864
rect 8895 833 8907 836
rect 8849 827 8907 833
rect 8938 756 8944 808
rect 8996 756 9002 808
rect 9048 805 9076 836
rect 9953 833 9965 867
rect 9999 864 10011 867
rect 13906 864 13912 876
rect 9999 836 10640 864
rect 9999 833 10011 836
rect 9953 827 10011 833
rect 10612 805 10640 836
rect 13372 836 13912 864
rect 13372 805 13400 836
rect 13906 824 13912 836
rect 13964 824 13970 876
rect 15841 867 15899 873
rect 15841 864 15853 867
rect 15672 836 15853 864
rect 15672 805 15700 836
rect 15841 833 15853 836
rect 15887 833 15899 867
rect 15841 827 15899 833
rect 17221 867 17279 873
rect 17221 833 17233 867
rect 17267 864 17279 867
rect 19797 867 19855 873
rect 17267 836 17448 864
rect 17267 833 17279 836
rect 17221 827 17279 833
rect 9033 799 9091 805
rect 9033 765 9045 799
rect 9079 765 9091 799
rect 9033 759 9091 765
rect 9125 799 9183 805
rect 9125 765 9137 799
rect 9171 796 9183 799
rect 9309 799 9367 805
rect 9309 796 9321 799
rect 9171 768 9321 796
rect 9171 765 9183 768
rect 9125 759 9183 765
rect 9309 765 9321 768
rect 9355 765 9367 799
rect 9309 759 9367 765
rect 9401 799 9459 805
rect 9401 765 9413 799
rect 9447 796 9459 799
rect 9585 799 9643 805
rect 9585 796 9597 799
rect 9447 768 9597 796
rect 9447 765 9459 768
rect 9401 759 9459 765
rect 9585 765 9597 768
rect 9631 765 9643 799
rect 9585 759 9643 765
rect 9677 799 9735 805
rect 9677 765 9689 799
rect 9723 796 9735 799
rect 9861 799 9919 805
rect 9861 796 9873 799
rect 9723 768 9873 796
rect 9723 765 9735 768
rect 9677 759 9735 765
rect 9861 765 9873 768
rect 9907 765 9919 799
rect 9861 759 9919 765
rect 10505 799 10563 805
rect 10505 765 10517 799
rect 10551 765 10563 799
rect 10505 759 10563 765
rect 10597 799 10655 805
rect 10597 765 10609 799
rect 10643 765 10655 799
rect 10597 759 10655 765
rect 13357 799 13415 805
rect 13357 765 13369 799
rect 13403 765 13415 799
rect 13357 759 13415 765
rect 13725 799 13783 805
rect 13725 765 13737 799
rect 13771 765 13783 799
rect 13725 759 13783 765
rect 13817 799 13875 805
rect 13817 765 13829 799
rect 13863 796 13875 799
rect 14001 799 14059 805
rect 14001 796 14013 799
rect 13863 768 14013 796
rect 13863 765 13875 768
rect 13817 759 13875 765
rect 14001 765 14013 768
rect 14047 765 14059 799
rect 14001 759 14059 765
rect 14093 799 14151 805
rect 14093 765 14105 799
rect 14139 796 14151 799
rect 14277 799 14335 805
rect 14277 796 14289 799
rect 14139 768 14289 796
rect 14139 765 14151 768
rect 14093 759 14151 765
rect 14277 765 14289 768
rect 14323 765 14335 799
rect 14277 759 14335 765
rect 14369 799 14427 805
rect 14369 765 14381 799
rect 14415 796 14427 799
rect 14553 799 14611 805
rect 14553 796 14565 799
rect 14415 768 14565 796
rect 14415 765 14427 768
rect 14369 759 14427 765
rect 14553 765 14565 768
rect 14599 765 14611 799
rect 14553 759 14611 765
rect 14645 799 14703 805
rect 14645 765 14657 799
rect 14691 796 14703 799
rect 14829 799 14887 805
rect 14829 796 14841 799
rect 14691 768 14841 796
rect 14691 765 14703 768
rect 14645 759 14703 765
rect 14829 765 14841 768
rect 14875 765 14887 799
rect 14829 759 14887 765
rect 14921 799 14979 805
rect 14921 765 14933 799
rect 14967 796 14979 799
rect 15105 799 15163 805
rect 15105 796 15117 799
rect 14967 768 15117 796
rect 14967 765 14979 768
rect 14921 759 14979 765
rect 15105 765 15117 768
rect 15151 765 15163 799
rect 15105 759 15163 765
rect 15657 799 15715 805
rect 15657 765 15669 799
rect 15703 765 15715 799
rect 15657 759 15715 765
rect 15749 799 15807 805
rect 15749 765 15761 799
rect 15795 765 15807 799
rect 15749 759 15807 765
rect 10520 728 10548 759
rect 10689 731 10747 737
rect 10689 728 10701 731
rect 10520 700 10701 728
rect 10689 697 10701 700
rect 10735 697 10747 731
rect 10689 691 10747 697
rect 13265 731 13323 737
rect 13265 697 13277 731
rect 13311 728 13323 731
rect 13740 728 13768 759
rect 13311 700 13768 728
rect 15197 731 15255 737
rect 13311 697 13323 700
rect 13265 691 13323 697
rect 15197 697 15209 731
rect 15243 728 15255 731
rect 15764 728 15792 759
rect 17310 756 17316 808
rect 17368 756 17374 808
rect 17420 805 17448 836
rect 19797 833 19809 867
rect 19843 864 19855 867
rect 19843 836 20116 864
rect 19843 833 19855 836
rect 19797 827 19855 833
rect 17405 799 17463 805
rect 17405 765 17417 799
rect 17451 765 17463 799
rect 17405 759 17463 765
rect 17497 799 17555 805
rect 17497 765 17509 799
rect 17543 796 17555 799
rect 17681 799 17739 805
rect 17681 796 17693 799
rect 17543 768 17693 796
rect 17543 765 17555 768
rect 17497 759 17555 765
rect 17681 765 17693 768
rect 17727 765 17739 799
rect 17681 759 17739 765
rect 17773 799 17831 805
rect 17773 765 17785 799
rect 17819 796 17831 799
rect 17957 799 18015 805
rect 17957 796 17969 799
rect 17819 768 17969 796
rect 17819 765 17831 768
rect 17773 759 17831 765
rect 17957 765 17969 768
rect 18003 765 18015 799
rect 17957 759 18015 765
rect 18049 799 18107 805
rect 18049 765 18061 799
rect 18095 796 18107 799
rect 18233 799 18291 805
rect 18233 796 18245 799
rect 18095 768 18245 796
rect 18095 765 18107 768
rect 18049 759 18107 765
rect 18233 765 18245 768
rect 18279 765 18291 799
rect 18233 759 18291 765
rect 18325 799 18383 805
rect 18325 765 18337 799
rect 18371 796 18383 799
rect 18693 799 18751 805
rect 18693 796 18705 799
rect 18371 768 18705 796
rect 18371 765 18383 768
rect 18325 759 18383 765
rect 18693 765 18705 768
rect 18739 765 18751 799
rect 18693 759 18751 765
rect 19886 756 19892 808
rect 19944 756 19950 808
rect 20088 805 20116 836
rect 20073 799 20131 805
rect 20073 765 20085 799
rect 20119 765 20131 799
rect 20073 759 20131 765
rect 20165 799 20223 805
rect 20165 765 20177 799
rect 20211 796 20223 799
rect 20349 799 20407 805
rect 20349 796 20361 799
rect 20211 768 20361 796
rect 20211 765 20223 768
rect 20165 759 20223 765
rect 20349 765 20361 768
rect 20395 765 20407 799
rect 20349 759 20407 765
rect 20441 799 20499 805
rect 20441 765 20453 799
rect 20487 796 20499 799
rect 20625 799 20683 805
rect 20625 796 20637 799
rect 20487 768 20637 796
rect 20487 765 20499 768
rect 20441 759 20499 765
rect 20625 765 20637 768
rect 20671 765 20683 799
rect 20625 759 20683 765
rect 20717 799 20775 805
rect 20717 765 20729 799
rect 20763 796 20775 799
rect 20901 799 20959 805
rect 20901 796 20913 799
rect 20763 768 20913 796
rect 20763 765 20775 768
rect 20717 759 20775 765
rect 20901 765 20913 768
rect 20947 765 20959 799
rect 20901 759 20959 765
rect 15243 700 15792 728
rect 15243 697 15255 700
rect 15197 691 15255 697
rect 552 570 31648 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31648 570
rect 552 496 31648 518
<< via1 >>
rect 19064 21836 19116 21888
rect 26424 21836 26476 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 11436 21734 11488 21786
rect 11500 21734 11552 21786
rect 11564 21734 11616 21786
rect 11628 21734 11680 21786
rect 11692 21734 11744 21786
rect 19210 21734 19262 21786
rect 19274 21734 19326 21786
rect 19338 21734 19390 21786
rect 19402 21734 19454 21786
rect 19466 21734 19518 21786
rect 26984 21734 27036 21786
rect 27048 21734 27100 21786
rect 27112 21734 27164 21786
rect 27176 21734 27228 21786
rect 27240 21734 27292 21786
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 7288 21675 7340 21684
rect 7288 21641 7297 21675
rect 7297 21641 7331 21675
rect 7331 21641 7340 21675
rect 7288 21632 7340 21641
rect 7840 21675 7892 21684
rect 7840 21641 7849 21675
rect 7849 21641 7883 21675
rect 7883 21641 7892 21675
rect 7840 21632 7892 21641
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 8944 21675 8996 21684
rect 8944 21641 8953 21675
rect 8953 21641 8987 21675
rect 8987 21641 8996 21675
rect 8944 21632 8996 21641
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 10048 21675 10100 21684
rect 10048 21641 10057 21675
rect 10057 21641 10091 21675
rect 10091 21641 10100 21675
rect 10048 21632 10100 21641
rect 10600 21675 10652 21684
rect 10600 21641 10609 21675
rect 10609 21641 10643 21675
rect 10643 21641 10652 21675
rect 10600 21632 10652 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11796 21632 11848 21684
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 15200 21632 15252 21684
rect 15660 21675 15712 21684
rect 15660 21641 15669 21675
rect 15669 21641 15703 21675
rect 15703 21641 15712 21675
rect 15660 21632 15712 21641
rect 16120 21675 16172 21684
rect 16120 21641 16129 21675
rect 16129 21641 16163 21675
rect 16163 21641 16172 21675
rect 16120 21632 16172 21641
rect 16764 21675 16816 21684
rect 16764 21641 16773 21675
rect 16773 21641 16807 21675
rect 16807 21641 16816 21675
rect 16764 21632 16816 21641
rect 16948 21675 17000 21684
rect 16948 21641 16957 21675
rect 16957 21641 16991 21675
rect 16991 21641 17000 21675
rect 16948 21632 17000 21641
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 18328 21675 18380 21684
rect 18328 21641 18337 21675
rect 18337 21641 18371 21675
rect 18371 21641 18380 21675
rect 18328 21632 18380 21641
rect 19064 21564 19116 21616
rect 19340 21564 19392 21616
rect 23204 21632 23256 21684
rect 26056 21632 26108 21684
rect 26424 21675 26476 21684
rect 26424 21641 26433 21675
rect 26433 21641 26467 21675
rect 26467 21641 26476 21675
rect 26424 21632 26476 21641
rect 16580 21471 16632 21480
rect 16580 21437 16589 21471
rect 16589 21437 16623 21471
rect 16623 21437 16632 21471
rect 16580 21428 16632 21437
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 18880 21428 18932 21480
rect 19800 21496 19852 21548
rect 20720 21496 20772 21548
rect 19708 21471 19760 21480
rect 19708 21437 19717 21471
rect 19717 21437 19751 21471
rect 19751 21437 19760 21471
rect 19708 21428 19760 21437
rect 20352 21471 20404 21480
rect 20352 21437 20361 21471
rect 20361 21437 20395 21471
rect 20395 21437 20404 21471
rect 20352 21428 20404 21437
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 22100 21428 22152 21480
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 22744 21471 22796 21480
rect 22744 21437 22753 21471
rect 22753 21437 22787 21471
rect 22787 21437 22796 21471
rect 22744 21428 22796 21437
rect 23204 21428 23256 21480
rect 21732 21335 21784 21344
rect 21732 21301 21741 21335
rect 21741 21301 21775 21335
rect 21775 21301 21784 21335
rect 21732 21292 21784 21301
rect 23296 21292 23348 21344
rect 23664 21292 23716 21344
rect 23848 21403 23900 21412
rect 23848 21369 23857 21403
rect 23857 21369 23891 21403
rect 23891 21369 23900 21403
rect 23848 21360 23900 21369
rect 24860 21428 24912 21480
rect 28172 21564 28224 21616
rect 26056 21428 26108 21480
rect 26332 21428 26384 21480
rect 27252 21471 27304 21480
rect 27252 21437 27261 21471
rect 27261 21437 27295 21471
rect 27295 21437 27304 21471
rect 27252 21428 27304 21437
rect 27528 21471 27580 21480
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 28632 21471 28684 21480
rect 28632 21437 28641 21471
rect 28641 21437 28675 21471
rect 28675 21437 28684 21471
rect 28632 21428 28684 21437
rect 29000 21471 29052 21480
rect 29000 21437 29009 21471
rect 29009 21437 29043 21471
rect 29043 21437 29052 21471
rect 29000 21428 29052 21437
rect 29460 21471 29512 21480
rect 29460 21437 29469 21471
rect 29469 21437 29503 21471
rect 29503 21437 29512 21471
rect 29460 21428 29512 21437
rect 29736 21471 29788 21480
rect 29736 21437 29745 21471
rect 29745 21437 29779 21471
rect 29779 21437 29788 21471
rect 29736 21428 29788 21437
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 25964 21403 26016 21412
rect 25964 21369 25973 21403
rect 25973 21369 26007 21403
rect 26007 21369 26016 21403
rect 25964 21360 26016 21369
rect 28080 21292 28132 21344
rect 29276 21292 29328 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 12096 21190 12148 21242
rect 12160 21190 12212 21242
rect 12224 21190 12276 21242
rect 12288 21190 12340 21242
rect 12352 21190 12404 21242
rect 19870 21190 19922 21242
rect 19934 21190 19986 21242
rect 19998 21190 20050 21242
rect 20062 21190 20114 21242
rect 20126 21190 20178 21242
rect 27644 21190 27696 21242
rect 27708 21190 27760 21242
rect 27772 21190 27824 21242
rect 27836 21190 27888 21242
rect 27900 21190 27952 21242
rect 16580 21088 16632 21140
rect 21088 21088 21140 21140
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 12348 20995 12400 21004
rect 12348 20961 12357 20995
rect 12357 20961 12391 20995
rect 12391 20961 12400 20995
rect 12348 20952 12400 20961
rect 19800 21020 19852 21072
rect 23848 21131 23900 21140
rect 23848 21097 23857 21131
rect 23857 21097 23891 21131
rect 23891 21097 23900 21131
rect 23848 21088 23900 21097
rect 25688 21088 25740 21140
rect 25964 21088 26016 21140
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 18880 20995 18932 21004
rect 18880 20961 18889 20995
rect 18889 20961 18923 20995
rect 18923 20961 18932 20995
rect 18880 20952 18932 20961
rect 19984 20995 20036 21004
rect 19984 20961 19993 20995
rect 19993 20961 20027 20995
rect 20027 20961 20036 20995
rect 19984 20952 20036 20961
rect 24216 21020 24268 21072
rect 28172 21088 28224 21140
rect 29000 21088 29052 21140
rect 29460 21088 29512 21140
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 23388 20995 23440 21004
rect 23388 20961 23397 20995
rect 23397 20961 23431 20995
rect 23431 20961 23440 20995
rect 23388 20952 23440 20961
rect 23480 20995 23532 21004
rect 23480 20961 23489 20995
rect 23489 20961 23523 20995
rect 23523 20961 23532 20995
rect 23480 20952 23532 20961
rect 24032 20995 24084 21004
rect 24032 20961 24041 20995
rect 24041 20961 24075 20995
rect 24075 20961 24084 20995
rect 24032 20952 24084 20961
rect 23664 20884 23716 20936
rect 24952 20995 25004 21004
rect 24952 20961 24961 20995
rect 24961 20961 24995 20995
rect 24995 20961 25004 20995
rect 24952 20952 25004 20961
rect 26240 20995 26292 21004
rect 26240 20961 26249 20995
rect 26249 20961 26283 20995
rect 26283 20961 26292 20995
rect 26240 20952 26292 20961
rect 28080 20952 28132 21004
rect 28816 20995 28868 21004
rect 28816 20961 28825 20995
rect 28825 20961 28859 20995
rect 28859 20961 28868 20995
rect 28816 20952 28868 20961
rect 29184 20995 29236 21004
rect 29184 20961 29193 20995
rect 29193 20961 29227 20995
rect 29227 20961 29236 20995
rect 29184 20952 29236 20961
rect 29276 20995 29328 21004
rect 29276 20961 29285 20995
rect 29285 20961 29319 20995
rect 29319 20961 29328 20995
rect 29276 20952 29328 20961
rect 23296 20816 23348 20868
rect 15016 20748 15068 20800
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 18512 20791 18564 20800
rect 18512 20757 18521 20791
rect 18521 20757 18555 20791
rect 18555 20757 18564 20791
rect 18512 20748 18564 20757
rect 20812 20748 20864 20800
rect 27436 20748 27488 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 11436 20646 11488 20698
rect 11500 20646 11552 20698
rect 11564 20646 11616 20698
rect 11628 20646 11680 20698
rect 11692 20646 11744 20698
rect 19210 20646 19262 20698
rect 19274 20646 19326 20698
rect 19338 20646 19390 20698
rect 19402 20646 19454 20698
rect 19466 20646 19518 20698
rect 26984 20646 27036 20698
rect 27048 20646 27100 20698
rect 27112 20646 27164 20698
rect 27176 20646 27228 20698
rect 27240 20646 27292 20698
rect 12348 20587 12400 20596
rect 12348 20553 12357 20587
rect 12357 20553 12391 20587
rect 12391 20553 12400 20587
rect 12348 20544 12400 20553
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 19984 20544 20036 20596
rect 23388 20544 23440 20596
rect 29184 20544 29236 20596
rect 1400 20340 1452 20392
rect 1124 20272 1176 20324
rect 3332 20340 3384 20392
rect 6460 20383 6512 20392
rect 6460 20349 6469 20383
rect 6469 20349 6503 20383
rect 6503 20349 6512 20383
rect 6460 20340 6512 20349
rect 11244 20383 11296 20392
rect 11244 20349 11253 20383
rect 11253 20349 11287 20383
rect 11287 20349 11296 20383
rect 11244 20340 11296 20349
rect 1216 20204 1268 20256
rect 1768 20204 1820 20256
rect 3700 20204 3752 20256
rect 8760 20204 8812 20256
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 16488 20383 16540 20392
rect 16488 20349 16497 20383
rect 16497 20349 16531 20383
rect 16531 20349 16540 20383
rect 16488 20340 16540 20349
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 18512 20383 18564 20392
rect 18512 20349 18521 20383
rect 18521 20349 18555 20383
rect 18555 20349 18564 20383
rect 18512 20340 18564 20349
rect 19708 20383 19760 20392
rect 19708 20349 19717 20383
rect 19717 20349 19751 20383
rect 19751 20349 19760 20383
rect 19708 20340 19760 20349
rect 20812 20383 20864 20392
rect 20812 20349 20821 20383
rect 20821 20349 20855 20383
rect 20855 20349 20864 20383
rect 20812 20340 20864 20349
rect 24400 20383 24452 20392
rect 24400 20349 24409 20383
rect 24409 20349 24443 20383
rect 24443 20349 24452 20383
rect 24400 20340 24452 20349
rect 27436 20383 27488 20392
rect 27436 20349 27445 20383
rect 27445 20349 27479 20383
rect 27479 20349 27488 20383
rect 27436 20340 27488 20349
rect 29000 20383 29052 20392
rect 29000 20349 29009 20383
rect 29009 20349 29043 20383
rect 29043 20349 29052 20383
rect 29000 20340 29052 20349
rect 14280 20204 14332 20256
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 19064 20204 19116 20256
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 26700 20247 26752 20256
rect 26700 20213 26709 20247
rect 26709 20213 26743 20247
rect 26743 20213 26752 20247
rect 26700 20204 26752 20213
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 12096 20102 12148 20154
rect 12160 20102 12212 20154
rect 12224 20102 12276 20154
rect 12288 20102 12340 20154
rect 12352 20102 12404 20154
rect 19870 20102 19922 20154
rect 19934 20102 19986 20154
rect 19998 20102 20050 20154
rect 20062 20102 20114 20154
rect 20126 20102 20178 20154
rect 27644 20102 27696 20154
rect 27708 20102 27760 20154
rect 27772 20102 27824 20154
rect 27836 20102 27888 20154
rect 27900 20102 27952 20154
rect 1124 20043 1176 20052
rect 1124 20009 1133 20043
rect 1133 20009 1167 20043
rect 1167 20009 1176 20043
rect 1124 20000 1176 20009
rect 1400 20043 1452 20052
rect 1400 20009 1409 20043
rect 1409 20009 1443 20043
rect 1443 20009 1452 20043
rect 1400 20000 1452 20009
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 6460 20043 6512 20052
rect 6460 20009 6469 20043
rect 6469 20009 6503 20043
rect 6503 20009 6512 20043
rect 6460 20000 6512 20009
rect 11244 20000 11296 20052
rect 17316 20000 17368 20052
rect 19708 20043 19760 20052
rect 19708 20009 19717 20043
rect 19717 20009 19751 20043
rect 19751 20009 19760 20043
rect 19708 20000 19760 20009
rect 24400 20000 24452 20052
rect 1216 19907 1268 19916
rect 1216 19873 1225 19907
rect 1225 19873 1259 19907
rect 1259 19873 1268 19907
rect 1216 19864 1268 19873
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 3700 19907 3752 19916
rect 3700 19873 3709 19907
rect 3709 19873 3743 19907
rect 3743 19873 3752 19907
rect 3700 19864 3752 19873
rect 4252 19907 4304 19916
rect 4252 19873 4261 19907
rect 4261 19873 4295 19907
rect 4295 19873 4304 19907
rect 4252 19864 4304 19873
rect 2872 19796 2924 19848
rect 8760 19907 8812 19916
rect 8760 19873 8769 19907
rect 8769 19873 8803 19907
rect 8803 19873 8812 19907
rect 8760 19864 8812 19873
rect 9588 19907 9640 19916
rect 9588 19873 9597 19907
rect 9597 19873 9631 19907
rect 9631 19873 9640 19907
rect 9588 19864 9640 19873
rect 10324 19907 10376 19916
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 5540 19728 5592 19780
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 19064 19907 19116 19916
rect 19064 19873 19073 19907
rect 19073 19873 19107 19907
rect 19107 19873 19116 19907
rect 19064 19864 19116 19873
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 21456 19907 21508 19916
rect 21456 19873 21465 19907
rect 21465 19873 21499 19907
rect 21499 19873 21508 19907
rect 21456 19864 21508 19873
rect 26056 19907 26108 19916
rect 26056 19873 26065 19907
rect 26065 19873 26099 19907
rect 26099 19873 26108 19907
rect 26056 19864 26108 19873
rect 27252 19907 27304 19916
rect 27252 19873 27261 19907
rect 27261 19873 27295 19907
rect 27295 19873 27304 19907
rect 27252 19864 27304 19873
rect 28356 19907 28408 19916
rect 28356 19873 28365 19907
rect 28365 19873 28399 19907
rect 28399 19873 28408 19907
rect 28356 19864 28408 19873
rect 2780 19660 2832 19712
rect 4344 19660 4396 19712
rect 5448 19660 5500 19712
rect 8392 19660 8444 19712
rect 9772 19660 9824 19712
rect 10508 19660 10560 19712
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 12992 19660 13044 19712
rect 15200 19703 15252 19712
rect 15200 19669 15209 19703
rect 15209 19669 15243 19703
rect 15243 19669 15252 19703
rect 15200 19660 15252 19669
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 22836 19660 22888 19712
rect 26516 19703 26568 19712
rect 26516 19669 26525 19703
rect 26525 19669 26559 19703
rect 26559 19669 26568 19703
rect 26516 19660 26568 19669
rect 29184 19660 29236 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 11436 19558 11488 19610
rect 11500 19558 11552 19610
rect 11564 19558 11616 19610
rect 11628 19558 11680 19610
rect 11692 19558 11744 19610
rect 19210 19558 19262 19610
rect 19274 19558 19326 19610
rect 19338 19558 19390 19610
rect 19402 19558 19454 19610
rect 19466 19558 19518 19610
rect 26984 19558 27036 19610
rect 27048 19558 27100 19610
rect 27112 19558 27164 19610
rect 27176 19558 27228 19610
rect 27240 19558 27292 19610
rect 1492 19456 1544 19508
rect 4252 19456 4304 19508
rect 9588 19456 9640 19508
rect 10324 19456 10376 19508
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 12716 19456 12768 19508
rect 17224 19456 17276 19508
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 26056 19456 26108 19508
rect 27344 19456 27396 19508
rect 28356 19456 28408 19508
rect 29000 19456 29052 19508
rect 1492 19295 1544 19304
rect 1492 19261 1501 19295
rect 1501 19261 1535 19295
rect 1535 19261 1544 19295
rect 1492 19252 1544 19261
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 2780 19252 2832 19261
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 3516 19252 3568 19304
rect 4344 19295 4396 19304
rect 4344 19261 4353 19295
rect 4353 19261 4387 19295
rect 4387 19261 4396 19295
rect 4344 19252 4396 19261
rect 5448 19295 5500 19304
rect 5448 19261 5457 19295
rect 5457 19261 5491 19295
rect 5491 19261 5500 19295
rect 5448 19252 5500 19261
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 12624 19320 12676 19372
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 18604 19320 18656 19372
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 3700 19116 3752 19168
rect 7288 19116 7340 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 14648 19116 14700 19168
rect 18788 19159 18840 19168
rect 18788 19125 18797 19159
rect 18797 19125 18831 19159
rect 18831 19125 18840 19159
rect 18788 19116 18840 19125
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 22836 19295 22888 19304
rect 22836 19261 22845 19295
rect 22845 19261 22879 19295
rect 22879 19261 22888 19295
rect 22836 19252 22888 19261
rect 26516 19252 26568 19304
rect 26700 19295 26752 19304
rect 26700 19261 26709 19295
rect 26709 19261 26743 19295
rect 26743 19261 26752 19295
rect 26700 19252 26752 19261
rect 27988 19252 28040 19304
rect 29184 19295 29236 19304
rect 29184 19261 29193 19295
rect 29193 19261 29227 19295
rect 29227 19261 29236 19295
rect 29184 19252 29236 19261
rect 23388 19116 23440 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 1492 18912 1544 18964
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 9312 18912 9364 18964
rect 17132 18912 17184 18964
rect 20812 18955 20864 18964
rect 20812 18921 20821 18955
rect 20821 18921 20855 18955
rect 20855 18921 20864 18955
rect 20812 18912 20864 18921
rect 27988 18955 28040 18964
rect 27988 18921 27997 18955
rect 27997 18921 28031 18955
rect 28031 18921 28040 18955
rect 27988 18912 28040 18921
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 3516 18776 3568 18828
rect 3700 18819 3752 18828
rect 3700 18785 3709 18819
rect 3709 18785 3743 18819
rect 3743 18785 3752 18819
rect 3700 18776 3752 18785
rect 7288 18819 7340 18828
rect 7288 18785 7297 18819
rect 7297 18785 7331 18819
rect 7331 18785 7340 18819
rect 7288 18776 7340 18785
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 12440 18844 12492 18896
rect 14648 18819 14700 18828
rect 14648 18785 14657 18819
rect 14657 18785 14691 18819
rect 14691 18785 14700 18819
rect 14648 18776 14700 18785
rect 16672 18776 16724 18828
rect 18788 18819 18840 18828
rect 18788 18785 18797 18819
rect 18797 18785 18831 18819
rect 18831 18785 18840 18819
rect 18788 18776 18840 18785
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 23388 18819 23440 18828
rect 23388 18785 23397 18819
rect 23397 18785 23431 18819
rect 23431 18785 23440 18819
rect 23388 18776 23440 18785
rect 28448 18819 28500 18828
rect 28448 18785 28457 18819
rect 28457 18785 28491 18819
rect 28491 18785 28500 18819
rect 28448 18776 28500 18785
rect 28724 18819 28776 18828
rect 28724 18785 28733 18819
rect 28733 18785 28767 18819
rect 28767 18785 28776 18819
rect 28724 18776 28776 18785
rect 6552 18572 6604 18624
rect 8024 18572 8076 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 14740 18572 14792 18624
rect 18880 18572 18932 18624
rect 25596 18572 25648 18624
rect 28540 18572 28592 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 1768 18368 1820 18420
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 9956 18368 10008 18420
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 21548 18368 21600 18420
rect 28448 18368 28500 18420
rect 28724 18411 28776 18420
rect 28724 18377 28733 18411
rect 28733 18377 28767 18411
rect 28767 18377 28776 18411
rect 28724 18368 28776 18377
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9680 18096 9732 18148
rect 5632 18028 5684 18080
rect 7472 18028 7524 18080
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 13544 18028 13596 18080
rect 14924 18071 14976 18080
rect 14924 18037 14933 18071
rect 14933 18037 14967 18071
rect 14967 18037 14976 18071
rect 14924 18028 14976 18037
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 19524 18207 19576 18216
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 18052 18028 18104 18080
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 19616 18028 19668 18080
rect 21824 18207 21876 18216
rect 21824 18173 21833 18207
rect 21833 18173 21867 18207
rect 21867 18173 21876 18207
rect 21824 18164 21876 18173
rect 25320 18164 25372 18216
rect 25596 18207 25648 18216
rect 25596 18173 25605 18207
rect 25605 18173 25639 18207
rect 25639 18173 25648 18207
rect 25596 18164 25648 18173
rect 28540 18164 28592 18216
rect 29736 18207 29788 18216
rect 29736 18173 29745 18207
rect 29745 18173 29779 18207
rect 29779 18173 29788 18207
rect 29736 18164 29788 18173
rect 24952 18028 25004 18080
rect 25780 18028 25832 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 1952 17824 2004 17876
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 19524 17824 19576 17876
rect 22100 17824 22152 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 29736 17824 29788 17876
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 4068 17731 4120 17740
rect 4068 17697 4077 17731
rect 4077 17697 4111 17731
rect 4111 17697 4120 17731
rect 4068 17688 4120 17697
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 9312 17731 9364 17740
rect 9312 17697 9321 17731
rect 9321 17697 9355 17731
rect 9355 17697 9364 17731
rect 9312 17688 9364 17697
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 18972 17731 19024 17740
rect 18972 17697 18981 17731
rect 18981 17697 19015 17731
rect 19015 17697 19024 17731
rect 18972 17688 19024 17697
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 23572 17731 23624 17740
rect 23572 17697 23581 17731
rect 23581 17697 23615 17731
rect 23615 17697 23624 17731
rect 23572 17688 23624 17697
rect 24952 17731 25004 17740
rect 24952 17697 24961 17731
rect 24961 17697 24995 17731
rect 24995 17697 25004 17731
rect 24952 17688 25004 17697
rect 25228 17731 25280 17740
rect 25228 17697 25237 17731
rect 25237 17697 25271 17731
rect 25271 17697 25280 17731
rect 25228 17688 25280 17697
rect 25780 17731 25832 17740
rect 25780 17697 25789 17731
rect 25789 17697 25823 17731
rect 25823 17697 25832 17731
rect 25780 17688 25832 17697
rect 27988 17688 28040 17740
rect 29552 17731 29604 17740
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 1308 17484 1360 17536
rect 7748 17484 7800 17536
rect 10048 17484 10100 17536
rect 12440 17484 12492 17536
rect 15016 17484 15068 17536
rect 20260 17484 20312 17536
rect 23020 17484 23072 17536
rect 26332 17484 26384 17536
rect 29000 17484 29052 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 1952 17280 2004 17332
rect 4068 17280 4120 17332
rect 9312 17280 9364 17332
rect 17592 17323 17644 17332
rect 17592 17289 17601 17323
rect 17601 17289 17635 17323
rect 17635 17289 17644 17323
rect 17592 17280 17644 17289
rect 23572 17280 23624 17332
rect 25228 17280 25280 17332
rect 29552 17280 29604 17332
rect 1308 17119 1360 17128
rect 1308 17085 1317 17119
rect 1317 17085 1351 17119
rect 1351 17085 1360 17119
rect 1308 17076 1360 17085
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5264 17076 5316 17128
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 13636 17076 13688 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 20260 17119 20312 17128
rect 20260 17085 20269 17119
rect 20269 17085 20303 17119
rect 20303 17085 20312 17119
rect 20260 17076 20312 17085
rect 23020 17119 23072 17128
rect 23020 17085 23029 17119
rect 23029 17085 23063 17119
rect 23063 17085 23072 17119
rect 23020 17076 23072 17085
rect 24216 17119 24268 17128
rect 24216 17085 24225 17119
rect 24225 17085 24259 17119
rect 24259 17085 24268 17119
rect 24216 17076 24268 17085
rect 26332 17119 26384 17128
rect 26332 17085 26341 17119
rect 26341 17085 26375 17119
rect 26375 17085 26384 17119
rect 26332 17076 26384 17085
rect 29000 17119 29052 17128
rect 29000 17085 29009 17119
rect 29009 17085 29043 17119
rect 29043 17085 29052 17119
rect 29000 17076 29052 17085
rect 30104 17119 30156 17128
rect 30104 17085 30113 17119
rect 30113 17085 30147 17119
rect 30147 17085 30156 17119
rect 30104 17076 30156 17085
rect 1768 16940 1820 16992
rect 8116 16940 8168 16992
rect 9772 16940 9824 16992
rect 11152 16940 11204 16992
rect 15384 16940 15436 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 20720 16940 20772 16992
rect 28080 16940 28132 16992
rect 29368 16940 29420 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 5264 16779 5316 16788
rect 5264 16745 5273 16779
rect 5273 16745 5307 16779
rect 5307 16745 5316 16779
rect 5264 16736 5316 16745
rect 9404 16736 9456 16788
rect 10784 16736 10836 16788
rect 13636 16779 13688 16788
rect 13636 16745 13645 16779
rect 13645 16745 13679 16779
rect 13679 16745 13688 16779
rect 13636 16736 13688 16745
rect 19248 16736 19300 16788
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10048 16600 10100 16609
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 15384 16643 15436 16652
rect 15384 16609 15393 16643
rect 15393 16609 15427 16643
rect 15427 16609 15436 16643
rect 15384 16600 15436 16609
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 18972 16643 19024 16652
rect 18972 16609 18981 16643
rect 18981 16609 19015 16643
rect 19015 16609 19024 16643
rect 18972 16600 19024 16609
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 27988 16779 28040 16788
rect 27988 16745 27997 16779
rect 27997 16745 28031 16779
rect 28031 16745 28040 16779
rect 27988 16736 28040 16745
rect 30104 16736 30156 16788
rect 30380 16668 30432 16720
rect 24952 16643 25004 16652
rect 24952 16609 24961 16643
rect 24961 16609 24995 16643
rect 24995 16609 25004 16643
rect 24952 16600 25004 16609
rect 26056 16643 26108 16652
rect 26056 16609 26065 16643
rect 26065 16609 26099 16643
rect 26099 16609 26108 16643
rect 26056 16600 26108 16609
rect 28080 16643 28132 16652
rect 28080 16609 28089 16643
rect 28089 16609 28123 16643
rect 28123 16609 28132 16643
rect 28080 16600 28132 16609
rect 29368 16643 29420 16652
rect 29368 16609 29377 16643
rect 29377 16609 29411 16643
rect 29411 16609 29420 16643
rect 29368 16600 29420 16609
rect 29920 16643 29972 16652
rect 29920 16609 29929 16643
rect 29929 16609 29963 16643
rect 29963 16609 29972 16643
rect 29920 16600 29972 16609
rect 7380 16396 7432 16448
rect 9588 16396 9640 16448
rect 15200 16439 15252 16448
rect 15200 16405 15209 16439
rect 15209 16405 15243 16439
rect 15243 16405 15252 16439
rect 15200 16396 15252 16405
rect 16948 16396 17000 16448
rect 22192 16396 22244 16448
rect 24124 16396 24176 16448
rect 25412 16439 25464 16448
rect 25412 16405 25421 16439
rect 25421 16405 25455 16439
rect 25455 16405 25464 16439
rect 25412 16396 25464 16405
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 4252 16192 4304 16244
rect 6092 16192 6144 16244
rect 13176 16192 13228 16244
rect 18972 16192 19024 16244
rect 24216 16235 24268 16244
rect 24216 16201 24225 16235
rect 24225 16201 24259 16235
rect 24259 16201 24268 16235
rect 24216 16192 24268 16201
rect 24952 16192 25004 16244
rect 26056 16192 26108 16244
rect 29920 16192 29972 16244
rect 4804 16056 4856 16108
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 15108 15988 15160 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 19248 16031 19300 16040
rect 19248 15997 19257 16031
rect 19257 15997 19291 16031
rect 19291 15997 19300 16031
rect 19248 15988 19300 15997
rect 22192 16031 22244 16040
rect 22192 15997 22201 16031
rect 22201 15997 22235 16031
rect 22235 15997 22244 16031
rect 22192 15988 22244 15997
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 25412 16031 25464 16040
rect 25412 15997 25421 16031
rect 25421 15997 25455 16031
rect 25455 15997 25464 16031
rect 25412 15988 25464 15997
rect 30104 16031 30156 16040
rect 30104 15997 30113 16031
rect 30113 15997 30147 16031
rect 30147 15997 30156 16031
rect 30104 15988 30156 15997
rect 30380 16031 30432 16040
rect 30380 15997 30389 16031
rect 30389 15997 30423 16031
rect 30423 15997 30432 16031
rect 30380 15988 30432 15997
rect 8944 15852 8996 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 11612 15852 11664 15904
rect 15752 15852 15804 15904
rect 17592 15852 17644 15904
rect 23112 15852 23164 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 4804 15648 4856 15700
rect 6552 15648 6604 15700
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 19248 15648 19300 15700
rect 30104 15691 30156 15700
rect 30104 15657 30113 15691
rect 30113 15657 30147 15691
rect 30147 15657 30156 15691
rect 30104 15648 30156 15657
rect 3976 15555 4028 15564
rect 3976 15521 3985 15555
rect 3985 15521 4019 15555
rect 4019 15521 4028 15555
rect 3976 15512 4028 15521
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 19616 15580 19668 15632
rect 22100 15555 22152 15564
rect 22100 15521 22109 15555
rect 22109 15521 22143 15555
rect 22143 15521 22152 15555
rect 22100 15512 22152 15521
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 29368 15555 29420 15564
rect 29368 15521 29377 15555
rect 29377 15521 29411 15555
rect 29411 15521 29420 15555
rect 29368 15512 29420 15521
rect 9312 15308 9364 15360
rect 14832 15308 14884 15360
rect 17224 15308 17276 15360
rect 22744 15308 22796 15360
rect 23664 15308 23716 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 4068 15104 4120 15156
rect 6276 15104 6328 15156
rect 19616 15147 19668 15156
rect 19616 15113 19625 15147
rect 19625 15113 19659 15147
rect 19659 15113 19668 15147
rect 19616 15104 19668 15113
rect 29368 15104 29420 15156
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 6460 14900 6512 14952
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 10416 14900 10468 14952
rect 11520 14900 11572 14952
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 18604 14900 18656 14952
rect 22744 14943 22796 14952
rect 22744 14909 22753 14943
rect 22753 14909 22787 14943
rect 22787 14909 22796 14943
rect 22744 14900 22796 14909
rect 23664 14943 23716 14952
rect 23664 14909 23673 14943
rect 23673 14909 23707 14943
rect 23707 14909 23716 14943
rect 23664 14900 23716 14909
rect 29000 14943 29052 14952
rect 29000 14909 29009 14943
rect 29009 14909 29043 14943
rect 29043 14909 29052 14943
rect 29000 14900 29052 14909
rect 31024 14900 31076 14952
rect 2780 14764 2832 14816
rect 9220 14764 9272 14816
rect 10876 14764 10928 14816
rect 11336 14764 11388 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 16396 14764 16448 14816
rect 20812 14764 20864 14816
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 30380 14764 30432 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 4160 14560 4212 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 22100 14603 22152 14612
rect 22100 14569 22109 14603
rect 22109 14569 22143 14603
rect 22143 14569 22152 14603
rect 22100 14560 22152 14569
rect 29000 14560 29052 14612
rect 31024 14603 31076 14612
rect 31024 14569 31033 14603
rect 31033 14569 31067 14603
rect 31067 14569 31076 14603
rect 31024 14560 31076 14569
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 20812 14467 20864 14476
rect 20812 14433 20821 14467
rect 20821 14433 20855 14467
rect 20855 14433 20864 14467
rect 20812 14424 20864 14433
rect 22468 14467 22520 14476
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 24124 14467 24176 14476
rect 24124 14433 24133 14467
rect 24133 14433 24167 14467
rect 24167 14433 24176 14467
rect 24124 14424 24176 14433
rect 30380 14467 30432 14476
rect 30380 14433 30389 14467
rect 30389 14433 30423 14467
rect 30423 14433 30432 14467
rect 30380 14424 30432 14433
rect 30840 14467 30892 14476
rect 30840 14433 30849 14467
rect 30849 14433 30883 14467
rect 30883 14433 30892 14467
rect 30840 14424 30892 14433
rect 2504 14220 2556 14272
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 16212 14220 16264 14272
rect 20260 14220 20312 14272
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 4160 14016 4212 14068
rect 10784 14016 10836 14068
rect 17592 14016 17644 14068
rect 22468 14016 22520 14068
rect 30840 14016 30892 14068
rect 19432 13948 19484 14000
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 10876 13855 10928 13864
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 22192 13855 22244 13864
rect 22192 13821 22201 13855
rect 22201 13821 22235 13855
rect 22235 13821 22244 13855
rect 22192 13812 22244 13821
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 30656 13855 30708 13864
rect 30656 13821 30665 13855
rect 30665 13821 30699 13855
rect 30699 13821 30708 13855
rect 30656 13812 30708 13821
rect 1952 13676 2004 13728
rect 6092 13676 6144 13728
rect 10968 13676 11020 13728
rect 11612 13676 11664 13728
rect 15292 13676 15344 13728
rect 29092 13719 29144 13728
rect 29092 13685 29101 13719
rect 29101 13685 29135 13719
rect 29135 13685 29144 13719
rect 29092 13676 29144 13685
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 3976 13472 4028 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 11796 13515 11848 13524
rect 11796 13481 11805 13515
rect 11805 13481 11839 13515
rect 11839 13481 11848 13515
rect 11796 13472 11848 13481
rect 17316 13472 17368 13524
rect 20996 13472 21048 13524
rect 22192 13472 22244 13524
rect 30656 13472 30708 13524
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 10968 13379 11020 13388
rect 10968 13345 10977 13379
rect 10977 13345 11011 13379
rect 11011 13345 11020 13379
rect 10968 13336 11020 13345
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 19432 13379 19484 13388
rect 19432 13345 19441 13379
rect 19441 13345 19475 13379
rect 19475 13345 19484 13379
rect 19432 13336 19484 13345
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 20260 13336 20312 13345
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 26148 13336 26200 13388
rect 26608 13379 26660 13388
rect 26608 13345 26617 13379
rect 26617 13345 26651 13379
rect 26651 13345 26660 13379
rect 26608 13336 26660 13345
rect 29092 13379 29144 13388
rect 29092 13345 29101 13379
rect 29101 13345 29135 13379
rect 29135 13345 29144 13379
rect 29092 13336 29144 13345
rect 30196 13379 30248 13388
rect 30196 13345 30205 13379
rect 30205 13345 30239 13379
rect 30239 13345 30248 13379
rect 30196 13336 30248 13345
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 7380 13132 7432 13184
rect 11980 13132 12032 13184
rect 15660 13132 15712 13184
rect 25320 13132 25372 13184
rect 26884 13132 26936 13184
rect 29000 13132 29052 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 4252 12928 4304 12980
rect 7012 12928 7064 12980
rect 13084 12928 13136 12980
rect 21548 12928 21600 12980
rect 26148 12971 26200 12980
rect 26148 12937 26157 12971
rect 26157 12937 26191 12971
rect 26191 12937 26200 12971
rect 26148 12928 26200 12937
rect 26608 12928 26660 12980
rect 30196 12928 30248 12980
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 6276 12724 6328 12776
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 13912 12656 13964 12708
rect 21824 12767 21876 12776
rect 21824 12733 21833 12767
rect 21833 12733 21867 12767
rect 21867 12733 21876 12767
rect 21824 12724 21876 12733
rect 25320 12767 25372 12776
rect 25320 12733 25329 12767
rect 25329 12733 25363 12767
rect 25363 12733 25372 12767
rect 25320 12724 25372 12733
rect 19432 12656 19484 12708
rect 26700 12767 26752 12776
rect 26700 12733 26709 12767
rect 26709 12733 26743 12767
rect 26743 12733 26752 12767
rect 26700 12724 26752 12733
rect 26884 12724 26936 12776
rect 29000 12767 29052 12776
rect 29000 12733 29009 12767
rect 29009 12733 29043 12767
rect 29043 12733 29052 12767
rect 29000 12724 29052 12733
rect 30840 12792 30892 12844
rect 2780 12588 2832 12640
rect 5632 12588 5684 12640
rect 11888 12588 11940 12640
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 20260 12588 20312 12640
rect 25044 12588 25096 12640
rect 28724 12588 28776 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 13912 12427 13964 12436
rect 13912 12393 13921 12427
rect 13921 12393 13955 12427
rect 13955 12393 13964 12427
rect 13912 12384 13964 12393
rect 19432 12384 19484 12436
rect 21824 12384 21876 12436
rect 26700 12384 26752 12436
rect 30840 12427 30892 12436
rect 30840 12393 30849 12427
rect 30849 12393 30883 12427
rect 30883 12393 30892 12427
rect 30840 12384 30892 12393
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 5632 12248 5684 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 15200 12248 15252 12300
rect 16304 12248 16356 12300
rect 20260 12291 20312 12300
rect 20260 12257 20269 12291
rect 20269 12257 20303 12291
rect 20303 12257 20312 12291
rect 20260 12248 20312 12257
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 26608 12291 26660 12300
rect 26608 12257 26617 12291
rect 26617 12257 26651 12291
rect 26651 12257 26660 12291
rect 26608 12248 26660 12257
rect 28724 12291 28776 12300
rect 28724 12257 28733 12291
rect 28733 12257 28767 12291
rect 28767 12257 28776 12291
rect 28724 12248 28776 12257
rect 30380 12291 30432 12300
rect 30380 12257 30389 12291
rect 30389 12257 30423 12291
rect 30423 12257 30432 12291
rect 30380 12248 30432 12257
rect 3240 12044 3292 12096
rect 6184 12044 6236 12096
rect 11336 12044 11388 12096
rect 15108 12044 15160 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 24952 12044 25004 12096
rect 28264 12087 28316 12096
rect 28264 12053 28273 12087
rect 28273 12053 28307 12087
rect 28307 12053 28316 12087
rect 28264 12044 28316 12053
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 13452 11840 13504 11892
rect 16304 11883 16356 11892
rect 16304 11849 16313 11883
rect 16313 11849 16347 11883
rect 16347 11849 16356 11883
rect 16304 11840 16356 11849
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 26608 11840 26660 11892
rect 30380 11883 30432 11892
rect 30380 11849 30389 11883
rect 30389 11849 30423 11883
rect 30423 11849 30432 11883
rect 30380 11840 30432 11849
rect 11336 11772 11388 11824
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6184 11636 6236 11645
rect 9680 11636 9732 11688
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 20444 11679 20496 11688
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 20444 11636 20496 11645
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 28264 11679 28316 11688
rect 28264 11645 28273 11679
rect 28273 11645 28307 11679
rect 28307 11645 28316 11679
rect 28264 11636 28316 11645
rect 30196 11679 30248 11688
rect 30196 11645 30205 11679
rect 30205 11645 30239 11679
rect 30239 11645 30248 11679
rect 30196 11636 30248 11645
rect 3516 11500 3568 11552
rect 11520 11500 11572 11552
rect 20904 11500 20956 11552
rect 28172 11500 28224 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 3516 11203 3568 11212
rect 3516 11169 3525 11203
rect 3525 11169 3559 11203
rect 3559 11169 3568 11203
rect 3516 11160 3568 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 13084 11296 13136 11348
rect 25872 11296 25924 11348
rect 30196 11296 30248 11348
rect 5632 11092 5684 11144
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 20628 11203 20680 11212
rect 20628 11169 20637 11203
rect 20637 11169 20671 11203
rect 20671 11169 20680 11203
rect 20628 11160 20680 11169
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 22836 11160 22888 11212
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 25964 11203 26016 11212
rect 25964 11169 25973 11203
rect 25973 11169 26007 11203
rect 26007 11169 26016 11203
rect 25964 11160 26016 11169
rect 28172 11203 28224 11212
rect 28172 11169 28181 11203
rect 28181 11169 28215 11203
rect 28215 11169 28224 11203
rect 28172 11160 28224 11169
rect 29368 11203 29420 11212
rect 29368 11169 29377 11203
rect 29377 11169 29411 11203
rect 29411 11169 29420 11203
rect 29368 11160 29420 11169
rect 16580 11024 16632 11076
rect 23848 11024 23900 11076
rect 4068 10956 4120 11008
rect 5908 10956 5960 11008
rect 8024 10956 8076 11008
rect 11796 10956 11848 11008
rect 14648 10956 14700 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 20720 10956 20772 11008
rect 26056 10956 26108 11008
rect 27344 10956 27396 11008
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 6000 10752 6052 10804
rect 10140 10752 10192 10804
rect 13728 10752 13780 10804
rect 16580 10795 16632 10804
rect 16580 10761 16589 10795
rect 16589 10761 16623 10795
rect 16623 10761 16632 10795
rect 16580 10752 16632 10761
rect 20628 10752 20680 10804
rect 25964 10752 26016 10804
rect 29368 10795 29420 10804
rect 29368 10761 29377 10795
rect 29377 10761 29411 10795
rect 29411 10761 29420 10795
rect 29368 10752 29420 10761
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 5908 10548 5960 10600
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 4068 10480 4120 10532
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 14648 10591 14700 10600
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 20720 10548 20772 10600
rect 21088 10591 21140 10600
rect 21088 10557 21097 10591
rect 21097 10557 21131 10591
rect 21131 10557 21140 10591
rect 21088 10548 21140 10557
rect 23848 10591 23900 10600
rect 23848 10557 23857 10591
rect 23857 10557 23891 10591
rect 23891 10557 23900 10591
rect 23848 10548 23900 10557
rect 24216 10548 24268 10600
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 26056 10591 26108 10600
rect 26056 10557 26065 10591
rect 26065 10557 26099 10591
rect 26099 10557 26108 10591
rect 26056 10548 26108 10557
rect 17960 10480 18012 10532
rect 27344 10591 27396 10600
rect 27344 10557 27353 10591
rect 27353 10557 27387 10591
rect 27387 10557 27396 10591
rect 27344 10548 27396 10557
rect 28816 10591 28868 10600
rect 28816 10557 28825 10591
rect 28825 10557 28859 10591
rect 28859 10557 28868 10591
rect 28816 10548 28868 10557
rect 3240 10412 3292 10464
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 17868 10412 17920 10464
rect 22928 10412 22980 10464
rect 23664 10412 23716 10464
rect 24768 10455 24820 10464
rect 24768 10421 24777 10455
rect 24777 10421 24811 10455
rect 24811 10421 24820 10455
rect 24768 10412 24820 10421
rect 25228 10412 25280 10464
rect 26700 10455 26752 10464
rect 26700 10421 26709 10455
rect 26709 10421 26743 10455
rect 26743 10421 26752 10455
rect 26700 10412 26752 10421
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 5172 10208 5224 10260
rect 3240 10115 3292 10124
rect 3240 10081 3249 10115
rect 3249 10081 3283 10115
rect 3283 10081 3292 10115
rect 3240 10072 3292 10081
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 3240 9868 3292 9920
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 9588 10208 9640 10260
rect 16764 10208 16816 10260
rect 21088 10208 21140 10260
rect 22836 10251 22888 10260
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 24216 10208 24268 10260
rect 24952 10208 25004 10260
rect 25136 10251 25188 10260
rect 25136 10217 25145 10251
rect 25145 10217 25179 10251
rect 25179 10217 25188 10251
rect 25136 10208 25188 10217
rect 28816 10251 28868 10260
rect 28816 10217 28825 10251
rect 28825 10217 28859 10251
rect 28859 10217 28868 10251
rect 28816 10208 28868 10217
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 19800 10115 19852 10124
rect 19800 10081 19809 10115
rect 19809 10081 19843 10115
rect 19843 10081 19852 10115
rect 19800 10072 19852 10081
rect 22928 10115 22980 10124
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 23664 10115 23716 10124
rect 23664 10081 23673 10115
rect 23673 10081 23707 10115
rect 23707 10081 23716 10115
rect 23664 10072 23716 10081
rect 24768 10140 24820 10192
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 26700 10115 26752 10124
rect 26700 10081 26709 10115
rect 26709 10081 26743 10115
rect 26743 10081 26752 10115
rect 26700 10072 26752 10081
rect 29552 10115 29604 10124
rect 29552 10081 29561 10115
rect 29561 10081 29595 10115
rect 29595 10081 29604 10115
rect 29552 10072 29604 10081
rect 7932 9868 7984 9920
rect 18420 9868 18472 9920
rect 26608 9868 26660 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 4896 9664 4948 9716
rect 16856 9664 16908 9716
rect 19800 9664 19852 9716
rect 29552 9664 29604 9716
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 4712 9460 4764 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 23204 9503 23256 9512
rect 23204 9469 23213 9503
rect 23213 9469 23247 9503
rect 23247 9469 23256 9503
rect 23204 9460 23256 9469
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 28816 9503 28868 9512
rect 28816 9469 28825 9503
rect 28825 9469 28859 9503
rect 28859 9469 28868 9503
rect 28816 9460 28868 9469
rect 3608 9324 3660 9376
rect 8576 9324 8628 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 15292 9324 15344 9376
rect 22652 9324 22704 9376
rect 26516 9324 26568 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 4712 9120 4764 9172
rect 8668 9163 8720 9172
rect 8668 9129 8677 9163
rect 8677 9129 8711 9163
rect 8711 9129 8720 9163
rect 8668 9120 8720 9129
rect 12808 9120 12860 9172
rect 17408 9120 17460 9172
rect 23204 9163 23256 9172
rect 23204 9129 23213 9163
rect 23213 9129 23247 9163
rect 23247 9129 23256 9163
rect 23204 9120 23256 9129
rect 28816 9163 28868 9172
rect 28816 9129 28825 9163
rect 28825 9129 28859 9163
rect 28859 9129 28868 9163
rect 28816 9120 28868 9129
rect 3608 9027 3660 9036
rect 3608 8993 3617 9027
rect 3617 8993 3651 9027
rect 3651 8993 3660 9027
rect 3608 8984 3660 8993
rect 7564 8984 7616 9036
rect 8576 9027 8628 9036
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 8576 8984 8628 8993
rect 11152 8984 11204 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 17868 9027 17920 9036
rect 17868 8993 17877 9027
rect 17877 8993 17911 9027
rect 17911 8993 17920 9027
rect 17868 8984 17920 8993
rect 19064 9027 19116 9036
rect 19064 8993 19073 9027
rect 19073 8993 19107 9027
rect 19107 8993 19116 9027
rect 19064 8984 19116 8993
rect 22376 9027 22428 9036
rect 22376 8993 22385 9027
rect 22385 8993 22419 9027
rect 22419 8993 22428 9027
rect 22376 8984 22428 8993
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 24492 9027 24544 9036
rect 24492 8993 24501 9027
rect 24501 8993 24535 9027
rect 24535 8993 24544 9027
rect 24492 8984 24544 8993
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 29552 9027 29604 9036
rect 29552 8993 29561 9027
rect 29561 8993 29595 9027
rect 29595 8993 29604 9027
rect 29552 8984 29604 8993
rect 8024 8780 8076 8832
rect 15108 8780 15160 8832
rect 18972 8823 19024 8832
rect 18972 8789 18981 8823
rect 18981 8789 19015 8823
rect 19015 8789 19024 8823
rect 18972 8780 19024 8789
rect 19616 8780 19668 8832
rect 21916 8780 21968 8832
rect 26700 8780 26752 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 11152 8576 11204 8628
rect 17868 8576 17920 8628
rect 19064 8576 19116 8628
rect 22376 8576 22428 8628
rect 24492 8576 24544 8628
rect 29552 8576 29604 8628
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 8484 8372 8536 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11336 8372 11388 8424
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 17040 8415 17092 8424
rect 17040 8381 17049 8415
rect 17049 8381 17083 8415
rect 17083 8381 17092 8415
rect 17040 8372 17092 8381
rect 19616 8440 19668 8492
rect 21916 8415 21968 8424
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 24492 8415 24544 8424
rect 24492 8381 24501 8415
rect 24501 8381 24535 8415
rect 24535 8381 24544 8415
rect 24492 8372 24544 8381
rect 26700 8415 26752 8424
rect 26700 8381 26709 8415
rect 26709 8381 26743 8415
rect 26743 8381 26752 8415
rect 26700 8372 26752 8381
rect 29276 8415 29328 8424
rect 29276 8381 29285 8415
rect 29285 8381 29319 8415
rect 29319 8381 29328 8415
rect 29276 8372 29328 8381
rect 7472 8236 7524 8288
rect 7748 8236 7800 8288
rect 8576 8279 8628 8288
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 9036 8236 9088 8288
rect 15384 8236 15436 8288
rect 29092 8279 29144 8288
rect 29092 8245 29101 8279
rect 29101 8245 29135 8279
rect 29135 8245 29144 8279
rect 29092 8236 29144 8245
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8668 8032 8720 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 17040 8032 17092 8084
rect 24492 8032 24544 8084
rect 29276 8032 29328 8084
rect 7380 7964 7432 8016
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8024 7939 8076 7948
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 11244 7896 11296 7948
rect 13544 7939 13596 7948
rect 13544 7905 13553 7939
rect 13553 7905 13587 7939
rect 13587 7905 13596 7939
rect 13544 7896 13596 7905
rect 8484 7828 8536 7880
rect 15384 7939 15436 7948
rect 15384 7905 15393 7939
rect 15393 7905 15427 7939
rect 15427 7905 15436 7939
rect 15384 7896 15436 7905
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23480 7939 23532 7948
rect 23480 7905 23489 7939
rect 23489 7905 23523 7939
rect 23523 7905 23532 7939
rect 23480 7896 23532 7905
rect 25964 7939 26016 7948
rect 25964 7905 25973 7939
rect 25973 7905 26007 7939
rect 26007 7905 26016 7939
rect 25964 7896 26016 7905
rect 29092 7939 29144 7948
rect 29092 7905 29101 7939
rect 29101 7905 29135 7939
rect 29135 7905 29144 7939
rect 29092 7896 29144 7905
rect 23020 7760 23072 7812
rect 7380 7692 7432 7744
rect 11336 7692 11388 7744
rect 15200 7692 15252 7744
rect 21916 7692 21968 7744
rect 22744 7692 22796 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 11244 7531 11296 7540
rect 11244 7497 11253 7531
rect 11253 7497 11287 7531
rect 11287 7497 11296 7531
rect 11244 7488 11296 7497
rect 13544 7488 13596 7540
rect 20352 7488 20404 7540
rect 22652 7488 22704 7540
rect 25964 7488 26016 7540
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 17224 7284 17276 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 19800 7327 19852 7336
rect 19800 7293 19809 7327
rect 19809 7293 19843 7327
rect 19843 7293 19852 7327
rect 19800 7284 19852 7293
rect 23480 7420 23532 7472
rect 21916 7327 21968 7336
rect 21916 7293 21925 7327
rect 21925 7293 21959 7327
rect 21959 7293 21968 7327
rect 21916 7284 21968 7293
rect 22744 7327 22796 7336
rect 22744 7293 22753 7327
rect 22753 7293 22787 7327
rect 22787 7293 22796 7327
rect 22744 7284 22796 7293
rect 23020 7327 23072 7336
rect 23020 7293 23029 7327
rect 23029 7293 23063 7327
rect 23063 7293 23072 7327
rect 23020 7284 23072 7293
rect 25780 7327 25832 7336
rect 25780 7293 25789 7327
rect 25789 7293 25823 7327
rect 25823 7293 25832 7327
rect 25780 7284 25832 7293
rect 7748 7148 7800 7200
rect 9956 7148 10008 7200
rect 15200 7148 15252 7200
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 18236 7148 18288 7200
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 7656 6944 7708 6996
rect 17224 6944 17276 6996
rect 19800 6987 19852 6996
rect 19800 6953 19809 6987
rect 19809 6953 19843 6987
rect 19843 6953 19852 6987
rect 19800 6944 19852 6953
rect 25780 6944 25832 6996
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14096 6740 14148 6792
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 17776 6851 17828 6860
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 18052 6808 18104 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 23480 6876 23532 6928
rect 26056 6851 26108 6860
rect 26056 6817 26065 6851
rect 26065 6817 26099 6851
rect 26099 6817 26108 6851
rect 26056 6808 26108 6817
rect 6460 6604 6512 6656
rect 10048 6604 10100 6656
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 21916 6647 21968 6656
rect 21916 6613 21925 6647
rect 21925 6613 21959 6647
rect 21959 6613 21968 6647
rect 21916 6604 21968 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 13452 6400 13504 6452
rect 15936 6400 15988 6452
rect 26056 6400 26108 6452
rect 6460 6239 6512 6248
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 8208 6196 8260 6248
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 13636 6239 13688 6248
rect 13636 6205 13645 6239
rect 13645 6205 13679 6239
rect 13679 6205 13688 6239
rect 13636 6196 13688 6205
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 10232 6060 10284 6112
rect 11796 6060 11848 6112
rect 12624 6060 12676 6112
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 26056 6239 26108 6248
rect 26056 6205 26065 6239
rect 26065 6205 26099 6239
rect 26099 6205 26108 6239
rect 26056 6196 26108 6205
rect 22008 6060 22060 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 11152 5856 11204 5908
rect 11704 5856 11756 5908
rect 16672 5856 16724 5908
rect 26056 5856 26108 5908
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 10232 5763 10284 5772
rect 10232 5729 10241 5763
rect 10241 5729 10275 5763
rect 10275 5729 10284 5763
rect 10232 5720 10284 5729
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 12624 5763 12676 5772
rect 12624 5729 12633 5763
rect 12633 5729 12667 5763
rect 12667 5729 12676 5763
rect 12624 5720 12676 5729
rect 16396 5763 16448 5772
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 19616 5720 19668 5772
rect 20444 5763 20496 5772
rect 20444 5729 20453 5763
rect 20453 5729 20487 5763
rect 20487 5729 20496 5763
rect 20444 5720 20496 5729
rect 20812 5720 20864 5772
rect 22008 5763 22060 5772
rect 22008 5729 22017 5763
rect 22017 5729 22051 5763
rect 22051 5729 22060 5763
rect 22008 5720 22060 5729
rect 24952 5763 25004 5772
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 6460 5516 6512 5568
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 17132 5516 17184 5568
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 20720 5516 20772 5568
rect 22468 5516 22520 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 9496 5312 9548 5364
rect 16396 5312 16448 5364
rect 19616 5312 19668 5364
rect 20812 5312 20864 5364
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 9496 5151 9548 5160
rect 9496 5117 9505 5151
rect 9505 5117 9539 5151
rect 9539 5117 9548 5151
rect 9496 5108 9548 5117
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 20444 5244 20496 5296
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 19708 5108 19760 5160
rect 20720 5176 20772 5228
rect 21272 5151 21324 5160
rect 21272 5117 21281 5151
rect 21281 5117 21315 5151
rect 21315 5117 21324 5151
rect 21272 5108 21324 5117
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24584 5040 24636 5092
rect 7012 4972 7064 5024
rect 14924 5015 14976 5024
rect 14924 4981 14933 5015
rect 14933 4981 14967 5015
rect 14967 4981 14976 5015
rect 14924 4972 14976 4981
rect 24492 4972 24544 5024
rect 25596 5015 25648 5024
rect 25596 4981 25605 5015
rect 25605 4981 25639 5015
rect 25639 4981 25648 5015
rect 25596 4972 25648 4981
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 9496 4768 9548 4820
rect 21272 4768 21324 4820
rect 24584 4768 24636 4820
rect 24952 4811 25004 4820
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 11888 4632 11940 4684
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 24492 4675 24544 4684
rect 24492 4641 24501 4675
rect 24501 4641 24535 4675
rect 24535 4641 24544 4675
rect 24492 4632 24544 4641
rect 25596 4632 25648 4684
rect 7012 4428 7064 4480
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 12072 4428 12124 4480
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 19616 4428 19668 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 8576 4224 8628 4276
rect 11888 4224 11940 4276
rect 17408 4224 17460 4276
rect 21824 4224 21876 4276
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 8300 4020 8352 4072
rect 24400 4088 24452 4140
rect 11428 4063 11480 4072
rect 11428 4029 11437 4063
rect 11437 4029 11471 4063
rect 11471 4029 11480 4063
rect 11428 4020 11480 4029
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 15660 4063 15712 4072
rect 15660 4029 15669 4063
rect 15669 4029 15703 4063
rect 15703 4029 15712 4063
rect 15660 4020 15712 4029
rect 17960 4063 18012 4072
rect 17960 4029 17969 4063
rect 17969 4029 18003 4063
rect 18003 4029 18012 4063
rect 17960 4020 18012 4029
rect 19616 4063 19668 4072
rect 19616 4029 19625 4063
rect 19625 4029 19659 4063
rect 19659 4029 19668 4063
rect 19616 4020 19668 4029
rect 25136 4020 25188 4072
rect 25780 4063 25832 4072
rect 25780 4029 25789 4063
rect 25789 4029 25823 4063
rect 25823 4029 25832 4063
rect 25780 4020 25832 4029
rect 26884 4063 26936 4072
rect 26884 4029 26893 4063
rect 26893 4029 26927 4063
rect 26927 4029 26936 4063
rect 26884 4020 26936 4029
rect 6736 3884 6788 3936
rect 10232 3884 10284 3936
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 20260 3884 20312 3936
rect 24492 3884 24544 3936
rect 25596 3927 25648 3936
rect 25596 3893 25605 3927
rect 25605 3893 25639 3927
rect 25639 3893 25648 3927
rect 25596 3884 25648 3893
rect 26148 3927 26200 3936
rect 26148 3893 26157 3927
rect 26157 3893 26191 3927
rect 26191 3893 26200 3927
rect 26148 3884 26200 3893
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 17960 3680 18012 3732
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 12624 3544 12676 3596
rect 12992 3544 13044 3596
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 25136 3680 25188 3732
rect 25780 3680 25832 3732
rect 26884 3680 26936 3732
rect 20260 3612 20312 3664
rect 24492 3587 24544 3596
rect 24492 3553 24501 3587
rect 24501 3553 24535 3587
rect 24535 3553 24544 3587
rect 24492 3544 24544 3553
rect 25596 3612 25648 3664
rect 26148 3544 26200 3596
rect 27528 3587 27580 3596
rect 27528 3553 27537 3587
rect 27537 3553 27571 3587
rect 27571 3553 27580 3587
rect 27528 3544 27580 3553
rect 6920 3340 6972 3392
rect 8668 3340 8720 3392
rect 12900 3340 12952 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 19708 3340 19760 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 8392 3136 8444 3188
rect 12624 3179 12676 3188
rect 12624 3145 12633 3179
rect 12633 3145 12667 3179
rect 12667 3145 12676 3179
rect 12624 3136 12676 3145
rect 12992 3179 13044 3188
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 18052 3136 18104 3188
rect 27528 3136 27580 3188
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 8668 2975 8720 2984
rect 8668 2941 8677 2975
rect 8677 2941 8711 2975
rect 8711 2941 8720 2975
rect 8668 2932 8720 2941
rect 11060 2975 11112 2984
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 19708 2975 19760 2984
rect 19708 2941 19717 2975
rect 19717 2941 19751 2975
rect 19751 2941 19760 2975
rect 19708 2932 19760 2941
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 26516 2975 26568 2984
rect 26516 2941 26525 2975
rect 26525 2941 26559 2975
rect 26559 2941 26568 2975
rect 26516 2932 26568 2941
rect 7564 2796 7616 2848
rect 11704 2796 11756 2848
rect 13728 2796 13780 2848
rect 13820 2796 13872 2848
rect 14280 2796 14332 2848
rect 18788 2796 18840 2848
rect 23940 2796 23992 2848
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 11060 2592 11112 2644
rect 11612 2592 11664 2644
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 11060 2456 11112 2508
rect 15844 2635 15896 2644
rect 15844 2601 15853 2635
rect 15853 2601 15887 2635
rect 15887 2601 15896 2635
rect 15844 2592 15896 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 26516 2592 26568 2644
rect 11244 2388 11296 2440
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 15568 2456 15620 2508
rect 18788 2499 18840 2508
rect 18788 2465 18797 2499
rect 18797 2465 18831 2499
rect 18831 2465 18840 2499
rect 18788 2456 18840 2465
rect 20628 2456 20680 2508
rect 23940 2499 23992 2508
rect 23940 2465 23949 2499
rect 23949 2465 23983 2499
rect 23983 2465 23992 2499
rect 23940 2456 23992 2465
rect 9036 2252 9088 2304
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 11060 2091 11112 2100
rect 11060 2057 11069 2091
rect 11069 2057 11103 2091
rect 11103 2057 11112 2091
rect 11060 2048 11112 2057
rect 11244 2048 11296 2100
rect 15568 2091 15620 2100
rect 15568 2057 15577 2091
rect 15577 2057 15611 2091
rect 15611 2057 15620 2091
rect 15568 2048 15620 2057
rect 20628 2091 20680 2100
rect 20628 2057 20637 2091
rect 20637 2057 20671 2091
rect 20671 2057 20680 2091
rect 20628 2048 20680 2057
rect 9036 1887 9088 1896
rect 9036 1853 9045 1887
rect 9045 1853 9079 1887
rect 9079 1853 9088 1887
rect 9036 1844 9088 1853
rect 10416 1912 10468 1964
rect 10876 1887 10928 1896
rect 10876 1853 10885 1887
rect 10885 1853 10919 1887
rect 10919 1853 10928 1887
rect 10876 1844 10928 1853
rect 13544 1887 13596 1896
rect 13544 1853 13553 1887
rect 13553 1853 13587 1887
rect 13587 1853 13596 1887
rect 13544 1844 13596 1853
rect 16304 1887 16356 1896
rect 16304 1853 16313 1887
rect 16313 1853 16347 1887
rect 16347 1853 16356 1887
rect 16304 1844 16356 1853
rect 21088 1912 21140 1964
rect 18604 1776 18656 1828
rect 8668 1751 8720 1760
rect 8668 1717 8677 1751
rect 8677 1717 8711 1751
rect 8711 1717 8720 1751
rect 8668 1708 8720 1717
rect 13176 1708 13228 1760
rect 17224 1708 17276 1760
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 10876 1504 10928 1556
rect 16304 1504 16356 1556
rect 8668 1411 8720 1420
rect 8668 1377 8677 1411
rect 8677 1377 8711 1411
rect 8711 1377 8720 1411
rect 8668 1368 8720 1377
rect 10232 1411 10284 1420
rect 10232 1377 10241 1411
rect 10241 1377 10275 1411
rect 10275 1377 10284 1411
rect 10232 1368 10284 1377
rect 13176 1411 13228 1420
rect 13176 1377 13185 1411
rect 13185 1377 13219 1411
rect 13219 1377 13228 1411
rect 13176 1368 13228 1377
rect 16396 1411 16448 1420
rect 16396 1377 16405 1411
rect 16405 1377 16439 1411
rect 16439 1377 16448 1411
rect 16396 1368 16448 1377
rect 17224 1411 17276 1420
rect 17224 1377 17233 1411
rect 17233 1377 17267 1411
rect 17267 1377 17276 1411
rect 17224 1368 17276 1377
rect 21088 1436 21140 1488
rect 18696 1411 18748 1420
rect 18696 1377 18705 1411
rect 18705 1377 18739 1411
rect 18739 1377 18748 1411
rect 18696 1368 18748 1377
rect 20720 1411 20772 1420
rect 20720 1377 20729 1411
rect 20729 1377 20763 1411
rect 20763 1377 20772 1411
rect 20720 1368 20772 1377
rect 8944 1164 8996 1216
rect 13912 1164 13964 1216
rect 17316 1164 17368 1216
rect 19892 1207 19944 1216
rect 19892 1173 19901 1207
rect 19901 1173 19935 1207
rect 19935 1173 19944 1207
rect 19892 1164 19944 1173
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 10232 960 10284 1012
rect 16396 960 16448 1012
rect 18696 960 18748 1012
rect 20720 960 20772 1012
rect 8944 799 8996 808
rect 8944 765 8953 799
rect 8953 765 8987 799
rect 8987 765 8996 799
rect 8944 756 8996 765
rect 13912 824 13964 876
rect 17316 799 17368 808
rect 17316 765 17325 799
rect 17325 765 17359 799
rect 17359 765 17368 799
rect 17316 756 17368 765
rect 19892 799 19944 808
rect 19892 765 19901 799
rect 19901 765 19935 799
rect 19935 765 19944 799
rect 19892 756 19944 765
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
<< metal2 >>
rect 28630 22128 28686 22137
rect 28630 22063 28686 22072
rect 11794 21992 11850 22001
rect 11794 21927 11850 21936
rect 12254 21992 12310 22001
rect 12254 21927 12310 21936
rect 19706 21992 19762 22001
rect 19706 21927 19762 21936
rect 20350 21992 20406 22001
rect 20350 21927 20406 21936
rect 22650 21992 22706 22001
rect 22650 21927 22706 21936
rect 27526 21992 27582 22001
rect 27526 21927 27582 21936
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 11436 21788 11744 21797
rect 11436 21786 11442 21788
rect 11498 21786 11522 21788
rect 11578 21786 11602 21788
rect 11658 21786 11682 21788
rect 11738 21786 11744 21788
rect 11498 21734 11500 21786
rect 11680 21734 11682 21786
rect 11436 21732 11442 21734
rect 11498 21732 11522 21734
rect 11578 21732 11602 21734
rect 11658 21732 11682 21734
rect 11738 21732 11744 21734
rect 6182 21720 6238 21729
rect 6182 21655 6184 21664
rect 6236 21655 6238 21664
rect 6734 21720 6790 21729
rect 6734 21655 6736 21664
rect 6184 21626 6236 21632
rect 6788 21655 6790 21664
rect 7286 21720 7342 21729
rect 7286 21655 7288 21664
rect 6736 21626 6788 21632
rect 7340 21655 7342 21664
rect 7838 21720 7894 21729
rect 7838 21655 7840 21664
rect 7288 21626 7340 21632
rect 7892 21655 7894 21664
rect 8390 21720 8446 21729
rect 8390 21655 8392 21664
rect 7840 21626 7892 21632
rect 8444 21655 8446 21664
rect 8942 21720 8998 21729
rect 8942 21655 8944 21664
rect 8392 21626 8444 21632
rect 8996 21655 8998 21664
rect 9494 21720 9550 21729
rect 9494 21655 9496 21664
rect 8944 21626 8996 21632
rect 9548 21655 9550 21664
rect 10046 21720 10102 21729
rect 10046 21655 10048 21664
rect 9496 21626 9548 21632
rect 10100 21655 10102 21664
rect 10598 21720 10654 21729
rect 10598 21655 10600 21664
rect 10048 21626 10100 21632
rect 10652 21655 10654 21664
rect 11150 21720 11206 21729
rect 11436 21723 11744 21732
rect 11808 21690 11836 21927
rect 12268 21690 12296 21927
rect 19064 21888 19116 21894
rect 16762 21856 16818 21865
rect 19064 21830 19116 21836
rect 16762 21791 16818 21800
rect 12806 21720 12862 21729
rect 11150 21655 11152 21664
rect 10600 21626 10652 21632
rect 11204 21655 11206 21664
rect 11796 21684 11848 21690
rect 11152 21626 11204 21632
rect 11796 21626 11848 21632
rect 12256 21684 12308 21690
rect 12806 21655 12808 21664
rect 12256 21626 12308 21632
rect 12860 21655 12862 21664
rect 13542 21720 13598 21729
rect 13542 21655 13544 21664
rect 12808 21626 12860 21632
rect 13596 21655 13598 21664
rect 13910 21720 13966 21729
rect 13910 21655 13912 21664
rect 13544 21626 13596 21632
rect 13964 21655 13966 21664
rect 14462 21720 14518 21729
rect 14462 21655 14464 21664
rect 13912 21626 13964 21632
rect 14516 21655 14518 21664
rect 15198 21720 15254 21729
rect 15198 21655 15200 21664
rect 14464 21626 14516 21632
rect 15252 21655 15254 21664
rect 15658 21720 15714 21729
rect 15658 21655 15660 21664
rect 15200 21626 15252 21632
rect 15712 21655 15714 21664
rect 16118 21720 16174 21729
rect 16776 21690 16804 21791
rect 16946 21720 17002 21729
rect 16118 21655 16120 21664
rect 15660 21626 15712 21632
rect 16172 21655 16174 21664
rect 16764 21684 16816 21690
rect 16120 21626 16172 21632
rect 16946 21655 16948 21664
rect 16764 21626 16816 21632
rect 17000 21655 17002 21664
rect 17590 21720 17646 21729
rect 17590 21655 17592 21664
rect 16948 21626 17000 21632
rect 17644 21655 17646 21664
rect 18326 21720 18382 21729
rect 18326 21655 18328 21664
rect 17592 21626 17644 21632
rect 18380 21655 18382 21664
rect 18328 21626 18380 21632
rect 19076 21622 19104 21830
rect 19210 21788 19518 21797
rect 19210 21786 19216 21788
rect 19272 21786 19296 21788
rect 19352 21786 19376 21788
rect 19432 21786 19456 21788
rect 19512 21786 19518 21788
rect 19272 21734 19274 21786
rect 19454 21734 19456 21786
rect 19210 21732 19216 21734
rect 19272 21732 19296 21734
rect 19352 21732 19376 21734
rect 19432 21732 19456 21734
rect 19512 21732 19518 21734
rect 19210 21723 19518 21732
rect 19064 21616 19116 21622
rect 19340 21616 19392 21622
rect 19064 21558 19116 21564
rect 19338 21584 19340 21593
rect 19392 21584 19394 21593
rect 19338 21519 19394 21528
rect 19720 21486 19748 21927
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 12096 21244 12404 21253
rect 12096 21242 12102 21244
rect 12158 21242 12182 21244
rect 12238 21242 12262 21244
rect 12318 21242 12342 21244
rect 12398 21242 12404 21244
rect 12158 21190 12160 21242
rect 12340 21190 12342 21242
rect 12096 21188 12102 21190
rect 12158 21188 12182 21190
rect 12238 21188 12262 21190
rect 12318 21188 12342 21190
rect 12398 21188 12404 21190
rect 12096 21179 12404 21188
rect 16592 21146 16620 21422
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 17420 21010 17448 21422
rect 18892 21010 18920 21422
rect 19812 21078 19840 21490
rect 20364 21486 20392 21927
rect 20718 21856 20774 21865
rect 20718 21791 20774 21800
rect 22098 21856 22154 21865
rect 22098 21791 22154 21800
rect 20732 21554 20760 21791
rect 21546 21584 21602 21593
rect 20720 21548 20772 21554
rect 21546 21519 21602 21528
rect 20720 21490 20772 21496
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 19870 21244 20178 21253
rect 19870 21242 19876 21244
rect 19932 21242 19956 21244
rect 20012 21242 20036 21244
rect 20092 21242 20116 21244
rect 20172 21242 20178 21244
rect 19932 21190 19934 21242
rect 20114 21190 20116 21242
rect 19870 21188 19876 21190
rect 19932 21188 19956 21190
rect 20012 21188 20036 21190
rect 20092 21188 20116 21190
rect 20172 21188 20178 21190
rect 19870 21179 20178 21188
rect 21100 21146 21128 21422
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 19800 21072 19852 21078
rect 19800 21014 19852 21020
rect 21560 21010 21588 21519
rect 22112 21486 22140 21791
rect 22664 21486 22692 21927
rect 26424 21888 26476 21894
rect 22742 21856 22798 21865
rect 22742 21791 22798 21800
rect 24858 21856 24914 21865
rect 26424 21830 26476 21836
rect 24858 21791 24914 21800
rect 22756 21486 22784 21791
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23216 21486 23244 21626
rect 23478 21584 23534 21593
rect 23478 21519 23534 21528
rect 24030 21584 24086 21593
rect 24030 21519 24086 21528
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 21744 21146 21772 21286
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 12348 21004 12400 21010
rect 12348 20946 12400 20952
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 11436 20700 11744 20709
rect 11436 20698 11442 20700
rect 11498 20698 11522 20700
rect 11578 20698 11602 20700
rect 11658 20698 11682 20700
rect 11738 20698 11744 20700
rect 11498 20646 11500 20698
rect 11680 20646 11682 20698
rect 11436 20644 11442 20646
rect 11498 20644 11522 20646
rect 11578 20644 11602 20646
rect 11658 20644 11682 20646
rect 11738 20644 11744 20646
rect 11436 20635 11744 20644
rect 12360 20602 12388 20946
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 15028 20398 15056 20742
rect 16500 20398 16528 20742
rect 17512 20602 17540 20946
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 18524 20398 18552 20742
rect 19210 20700 19518 20709
rect 19210 20698 19216 20700
rect 19272 20698 19296 20700
rect 19352 20698 19376 20700
rect 19432 20698 19456 20700
rect 19512 20698 19518 20700
rect 19272 20646 19274 20698
rect 19454 20646 19456 20698
rect 19210 20644 19216 20646
rect 19272 20644 19296 20646
rect 19352 20644 19376 20646
rect 19432 20644 19456 20646
rect 19512 20644 19518 20646
rect 19210 20635 19518 20644
rect 19996 20602 20024 20946
rect 23308 20874 23336 21286
rect 23492 21010 23520 21519
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20824 20398 20852 20742
rect 23400 20602 23428 20946
rect 23676 20942 23704 21286
rect 23860 21146 23888 21354
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24044 21010 24072 21519
rect 24872 21486 24900 21791
rect 26436 21690 26464 21830
rect 26984 21788 27292 21797
rect 26984 21786 26990 21788
rect 27046 21786 27070 21788
rect 27126 21786 27150 21788
rect 27206 21786 27230 21788
rect 27286 21786 27292 21788
rect 27046 21734 27048 21786
rect 27228 21734 27230 21786
rect 26984 21732 26990 21734
rect 27046 21732 27070 21734
rect 27126 21732 27150 21734
rect 27206 21732 27230 21734
rect 27286 21732 27292 21734
rect 26984 21723 27292 21732
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 24950 21584 25006 21593
rect 24950 21519 25006 21528
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 21078 24256 21286
rect 24216 21072 24268 21078
rect 24216 21014 24268 21020
rect 24964 21010 24992 21519
rect 26068 21486 26096 21626
rect 27250 21584 27306 21593
rect 27250 21519 27306 21528
rect 27264 21486 27292 21519
rect 27540 21486 27568 21927
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 25964 21412 26016 21418
rect 25964 21354 26016 21360
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25700 21146 25728 21286
rect 25976 21146 26004 21354
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 1124 20324 1176 20330
rect 1124 20266 1176 20272
rect 1136 20058 1164 20266
rect 1216 20256 1268 20262
rect 1216 20198 1268 20204
rect 1124 20052 1176 20058
rect 1124 19994 1176 20000
rect 1228 19922 1256 20198
rect 1412 20058 1440 20334
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1780 19922 1808 20198
rect 3344 20058 3372 20334
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3712 19922 3740 20198
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 6472 20058 6500 20334
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 8772 19922 8800 20198
rect 11256 20058 11284 20334
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 12096 20156 12404 20165
rect 12096 20154 12102 20156
rect 12158 20154 12182 20156
rect 12238 20154 12262 20156
rect 12318 20154 12342 20156
rect 12398 20154 12404 20156
rect 12158 20102 12160 20154
rect 12340 20102 12342 20154
rect 12096 20100 12102 20102
rect 12158 20100 12182 20102
rect 12238 20100 12262 20102
rect 12318 20100 12342 20102
rect 12398 20100 12404 20102
rect 12096 20091 12404 20100
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 14292 19922 14320 20198
rect 16132 19922 16160 20198
rect 17328 20058 17356 20334
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 19076 19922 19104 20198
rect 19720 20058 19748 20334
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 19870 20156 20178 20165
rect 19870 20154 19876 20156
rect 19932 20154 19956 20156
rect 20012 20154 20036 20156
rect 20092 20154 20116 20156
rect 20172 20154 20178 20156
rect 19932 20102 19934 20154
rect 20114 20102 20116 20154
rect 19870 20100 19876 20102
rect 19932 20100 19956 20102
rect 20012 20100 20036 20102
rect 20092 20100 20116 20102
rect 20172 20100 20178 20102
rect 19870 20091 20178 20100
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 21468 19922 21496 20198
rect 24412 20058 24440 20334
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 1504 19514 1532 19858
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 2792 19310 2820 19654
rect 2884 19310 2912 19790
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 4264 19514 4292 19858
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4356 19310 4384 19654
rect 5460 19310 5488 19654
rect 5552 19310 5580 19722
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19310 8432 19654
rect 9600 19514 9628 19858
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9784 19310 9812 19654
rect 10336 19514 10364 19858
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10520 19310 10548 19654
rect 10612 19514 10640 19858
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 11436 19612 11744 19621
rect 11436 19610 11442 19612
rect 11498 19610 11522 19612
rect 11578 19610 11602 19612
rect 11658 19610 11682 19612
rect 11738 19610 11744 19612
rect 11498 19558 11500 19610
rect 11680 19558 11682 19610
rect 11436 19556 11442 19558
rect 11498 19556 11522 19558
rect 11578 19556 11602 19558
rect 11658 19556 11682 19558
rect 11738 19556 11744 19558
rect 11436 19547 11744 19556
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 12636 19378 12664 19654
rect 12728 19514 12756 19858
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 13004 19310 13032 19654
rect 15212 19310 15240 19654
rect 17236 19514 17264 19858
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 18616 19378 18644 19654
rect 19210 19612 19518 19621
rect 19210 19610 19216 19612
rect 19272 19610 19296 19612
rect 19352 19610 19376 19612
rect 19432 19610 19456 19612
rect 19512 19610 19518 19612
rect 19272 19558 19274 19610
rect 19454 19558 19456 19610
rect 19210 19556 19216 19558
rect 19272 19556 19296 19558
rect 19352 19556 19376 19558
rect 19432 19556 19456 19558
rect 19512 19556 19518 19558
rect 19210 19547 19518 19556
rect 20180 19514 20208 19858
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 22848 19310 22876 19654
rect 26068 19514 26096 19858
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26252 19417 26280 20946
rect 26344 19553 26372 21422
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27644 21244 27952 21253
rect 27644 21242 27650 21244
rect 27706 21242 27730 21244
rect 27786 21242 27810 21244
rect 27866 21242 27890 21244
rect 27946 21242 27952 21244
rect 27706 21190 27708 21242
rect 27888 21190 27890 21242
rect 27644 21188 27650 21190
rect 27706 21188 27730 21190
rect 27786 21188 27810 21190
rect 27866 21188 27890 21190
rect 27946 21188 27952 21190
rect 27644 21179 27952 21188
rect 28092 21010 28120 21286
rect 28184 21146 28212 21558
rect 28644 21486 28672 22063
rect 29734 21856 29790 21865
rect 29734 21791 29790 21800
rect 28814 21584 28870 21593
rect 28814 21519 28870 21528
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28828 21010 28856 21519
rect 29748 21486 29776 21791
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 29012 21146 29040 21422
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 29288 21010 29316 21286
rect 29472 21146 29500 21422
rect 29460 21140 29512 21146
rect 29460 21082 29512 21088
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 28816 21004 28868 21010
rect 28816 20946 28868 20952
rect 29184 21004 29236 21010
rect 29184 20946 29236 20952
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 26984 20700 27292 20709
rect 26984 20698 26990 20700
rect 27046 20698 27070 20700
rect 27126 20698 27150 20700
rect 27206 20698 27230 20700
rect 27286 20698 27292 20700
rect 27046 20646 27048 20698
rect 27228 20646 27230 20698
rect 26984 20644 26990 20646
rect 27046 20644 27070 20646
rect 27126 20644 27150 20646
rect 27206 20644 27230 20646
rect 27286 20644 27292 20646
rect 26984 20635 27292 20644
rect 27448 20398 27476 20742
rect 29196 20602 29224 20946
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 26700 20256 26752 20262
rect 26700 20198 26752 20204
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26330 19544 26386 19553
rect 26330 19479 26386 19488
rect 26238 19408 26294 19417
rect 26238 19343 26294 19352
rect 26528 19310 26556 19654
rect 26712 19310 26740 20198
rect 27644 20156 27952 20165
rect 27644 20154 27650 20156
rect 27706 20154 27730 20156
rect 27786 20154 27810 20156
rect 27866 20154 27890 20156
rect 27946 20154 27952 20156
rect 27706 20102 27708 20154
rect 27888 20102 27890 20154
rect 27644 20100 27650 20102
rect 27706 20100 27730 20102
rect 27786 20100 27810 20102
rect 27866 20100 27890 20102
rect 27946 20100 27952 20102
rect 27644 20091 27952 20100
rect 27252 19916 27304 19922
rect 28356 19916 28408 19922
rect 27304 19876 27384 19904
rect 27252 19858 27304 19864
rect 26984 19612 27292 19621
rect 26984 19610 26990 19612
rect 27046 19610 27070 19612
rect 27126 19610 27150 19612
rect 27206 19610 27230 19612
rect 27286 19610 27292 19612
rect 27046 19558 27048 19610
rect 27228 19558 27230 19610
rect 26984 19556 26990 19558
rect 27046 19556 27070 19558
rect 27126 19556 27150 19558
rect 27206 19556 27230 19558
rect 27286 19556 27292 19558
rect 26984 19547 27292 19556
rect 27356 19514 27384 19876
rect 28356 19858 28408 19864
rect 28368 19514 28396 19858
rect 29012 19514 29040 20334
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 29196 19310 29224 19654
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 1504 18970 1532 19246
rect 3528 18970 3556 19246
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3712 18834 3740 19110
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 7300 18834 7328 19110
rect 9324 18970 9352 19246
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 12452 18902 12480 19110
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 14660 18834 14688 19110
rect 17144 18970 17172 19246
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 18800 18834 18828 19110
rect 19870 19068 20178 19077
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 20824 18970 20852 19246
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 23400 18834 23428 19110
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 28000 18970 28028 19246
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 1780 18426 1808 18770
rect 3528 18426 3556 18770
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 6564 18222 6592 18566
rect 8036 18222 8064 18566
rect 9968 18426 9996 18770
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 12728 18222 12756 18566
rect 14752 18222 14780 18566
rect 16684 18426 16712 18770
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 18892 18222 18920 18566
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 21560 18426 21588 18770
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 25608 18222 25636 18566
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 28460 18426 28488 18770
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28552 18222 28580 18566
rect 28736 18426 28764 18770
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 21824 18216 21876 18222
rect 25320 18216 25372 18222
rect 21876 18164 22140 18170
rect 21824 18158 22140 18164
rect 25320 18158 25372 18164
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 1964 17882 1992 18158
rect 3896 17882 3924 18158
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 5644 17746 5672 18022
rect 7484 17746 7512 18022
rect 9692 17882 9720 18090
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 13556 17746 13584 18022
rect 14936 17746 14964 18022
rect 18064 17882 18092 18022
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18984 17746 19012 18022
rect 19536 17882 19564 18158
rect 21836 18142 22140 18158
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19628 17746 19656 18022
rect 19870 17980 20178 17989
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 22112 17882 22140 18142
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 24964 17746 24992 18022
rect 25332 17882 25360 18158
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25792 17746 25820 18022
rect 27644 17980 27952 17989
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 29748 17882 29776 18158
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 1308 17536 1360 17542
rect 1308 17478 1360 17484
rect 1320 17134 1348 17478
rect 1308 17128 1360 17134
rect 1308 17070 1360 17076
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16658 1808 16934
rect 1872 16794 1900 17682
rect 1964 17338 1992 17682
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4080 17338 4108 17682
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 7760 17134 7788 17478
rect 9324 17338 9352 17682
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4908 16794 4936 17070
rect 5276 16794 5304 17070
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 8128 16658 8156 16934
rect 9416 16794 9444 17070
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9784 16658 9812 16934
rect 10060 16658 10088 17478
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 12452 17134 12480 17478
rect 15028 17134 15056 17478
rect 17604 17338 17632 17682
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 20272 17134 20300 17478
rect 23032 17134 23060 17478
rect 23584 17338 23612 17682
rect 25240 17338 25268 17682
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 26344 17134 26372 17478
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 10796 16794 10824 17070
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 11164 16658 11192 16934
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 13648 16794 13676 17070
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 15396 16658 15424 16934
rect 16684 16658 16712 16934
rect 19260 16794 19288 17070
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 20732 16658 20760 16934
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4264 16250 4292 16594
rect 6104 16250 6132 16594
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4816 15706 4844 16050
rect 7392 16046 7420 16390
rect 9600 16046 9628 16390
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 13188 16250 13216 16594
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 15108 16040 15160 16046
rect 15212 16028 15240 16390
rect 16960 16046 16988 16390
rect 18984 16250 19012 16594
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 22204 16046 22232 16390
rect 24136 16046 24164 16390
rect 24228 16250 24256 17070
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 28000 16794 28028 17682
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17134 29040 17478
rect 29564 17338 29592 17682
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 28092 16658 28120 16934
rect 29380 16658 29408 16934
rect 30116 16794 30144 17070
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30380 16720 30432 16726
rect 30380 16662 30432 16668
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29920 16652 29972 16658
rect 29920 16594 29972 16600
rect 24964 16250 24992 16594
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 25424 16046 25452 16390
rect 26068 16250 26096 16594
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 29932 16250 29960 16594
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 30392 16046 30420 16662
rect 15160 16000 15240 16028
rect 16948 16040 17000 16046
rect 15108 15982 15160 15988
rect 16948 15982 17000 15988
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 6564 15706 6592 15982
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 8956 15570 8984 15846
rect 9416 15570 9444 15846
rect 11072 15706 11100 15982
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11624 15570 11652 15846
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 13188 15706 13216 15982
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 15764 15570 15792 15846
rect 17604 15570 17632 15846
rect 19260 15706 19288 15982
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 19870 15804 20178 15813
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 3988 15450 4016 15506
rect 3988 15422 4108 15450
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4080 15162 4108 15422
rect 6288 15162 6316 15506
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 9324 14958 9352 15302
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 14844 14958 14872 15302
rect 17236 14958 17264 15302
rect 19210 15260 19518 15269
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 19628 15162 19656 15574
rect 23124 15570 23152 15846
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 30116 15706 30144 15982
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14482 2820 14758
rect 4172 14618 4200 14894
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 6472 14618 6500 14894
rect 7668 14618 7696 14894
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 9232 14482 9260 14758
rect 10428 14618 10456 14894
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13870 2544 14214
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 4172 14074 4200 14418
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 6104 13818 6132 14418
rect 10796 14074 10824 14418
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10888 13870 10916 14758
rect 11348 14482 11376 14758
rect 11532 14618 11560 14894
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 14384 14482 14412 14758
rect 16408 14482 16436 14758
rect 18616 14618 18644 14894
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 20824 14482 20852 14758
rect 22112 14618 22140 15506
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 22756 14958 22784 15302
rect 23676 14958 23704 15302
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 29380 15162 29408 15506
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 24136 14482 24164 14758
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 29012 14618 29040 14894
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 30392 14482 30420 14758
rect 31036 14618 31064 14894
rect 31024 14612 31076 14618
rect 31024 14554 31076 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 11256 13870 11284 14214
rect 11436 14172 11744 14181
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11436 14107 11744 14116
rect 16224 13870 16252 14214
rect 17604 14074 17632 14418
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 6644 13864 6696 13870
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13394 1992 13670
rect 3988 13530 4016 13806
rect 6104 13790 6224 13818
rect 6644 13806 6696 13812
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 6104 13394 6132 13670
rect 6196 13530 6224 13790
rect 6656 13530 6684 13806
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 10980 13394 11008 13670
rect 11624 13394 11652 13670
rect 11808 13530 11836 13806
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 15304 13394 15332 13670
rect 17328 13530 17356 13806
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 19444 13394 19472 13942
rect 19870 13628 20178 13637
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 20272 13394 20300 14214
rect 22480 14074 22508 14418
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 25148 13870 25176 14214
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 30852 14074 30880 14418
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 30656 13864 30708 13870
rect 30656 13806 30708 13812
rect 21008 13530 21036 13806
rect 22204 13530 22232 13806
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 29104 13394 29132 13670
rect 30668 13530 30696 13806
rect 30656 13524 30708 13530
rect 30656 13466 30708 13472
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12782 2452 13126
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 4264 12986 4292 13330
rect 7024 12986 7052 13330
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7392 12782 7420 13126
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 11992 12782 12020 13126
rect 13096 12986 13124 13330
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 15672 12782 15700 13126
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 21560 12986 21588 13330
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 25332 12782 25360 13126
rect 26160 12986 26188 13330
rect 26620 12986 26648 13330
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26896 12782 26924 13126
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 29012 12782 29040 13126
rect 30208 12986 30236 13330
rect 30196 12980 30248 12986
rect 30196 12922 30248 12928
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26884 12776 26936 12782
rect 26884 12718 26936 12724
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12306 2820 12582
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 5000 12442 5028 12718
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5644 12306 5672 12582
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 3252 11694 3280 12038
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 6196 11694 6224 12038
rect 6288 11898 6316 12718
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12306 11928 12582
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 13924 12442 13952 12650
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 15212 12306 15240 12582
rect 19444 12442 19472 12650
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 20272 12306 20300 12582
rect 21836 12442 21864 12718
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 25056 12306 25084 12582
rect 26712 12442 26740 12718
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 28736 12306 28764 12582
rect 30852 12442 30880 12786
rect 30840 12436 30892 12442
rect 30840 12378 30892 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 28724 12300 28776 12306
rect 28724 12242 28776 12248
rect 30380 12300 30432 12306
rect 30380 12242 30432 12248
rect 9692 11898 9720 12242
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 11348 11830 11376 12038
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 13464 11898 13492 12242
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 15120 11694 15148 12038
rect 16316 11898 16344 12242
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 20456 11694 20484 12038
rect 22296 11898 22324 12242
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 24964 11694 24992 12038
rect 26620 11898 26648 12242
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 28276 11694 28304 12038
rect 30392 11898 30420 12242
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 28264 11688 28316 11694
rect 28264 11630 28316 11636
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 9692 11354 9720 11630
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 11532 11218 11560 11494
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 12096 11387 12404 11396
rect 13096 11354 13124 11630
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 20916 11218 20944 11494
rect 25884 11354 25912 11630
rect 28172 11552 28224 11558
rect 28172 11494 28224 11500
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 28184 11218 28212 11494
rect 30208 11354 30236 11630
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 4080 10538 4108 10950
rect 5644 10810 5672 11086
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5920 10606 5948 10950
rect 6012 10810 6040 11154
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 8036 10606 8064 10950
rect 10152 10810 10180 11154
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11436 10843 11744 10852
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 11808 10606 11836 10950
rect 13740 10810 13768 11154
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 14660 10606 14688 10950
rect 16592 10810 16620 11018
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10130 3280 10406
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 5184 10266 5212 10542
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 7668 10130 7696 10406
rect 9600 10266 9628 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9784 10130 9812 10406
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 16776 10266 16804 10542
rect 17972 10538 18000 10950
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 20640 10810 20668 11154
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20732 10606 20760 10950
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 17880 10130 17908 10406
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 21100 10266 21128 10542
rect 22848 10266 22876 11154
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 10606 23888 11018
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22940 10130 22968 10406
rect 23676 10130 23704 10406
rect 24228 10266 24256 10542
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24780 10198 24808 10406
rect 24964 10266 24992 10542
rect 25148 10266 25176 11154
rect 25976 10810 26004 11154
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 26068 10606 26096 10950
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 27356 10606 27384 10950
rect 29380 10810 29408 11154
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 26056 10600 26108 10606
rect 26056 10542 26108 10548
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 25240 10130 25268 10406
rect 26712 10130 26740 10406
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 28828 10266 28856 10542
rect 28816 10260 28868 10266
rect 28816 10202 28868 10208
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9518 3280 9862
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4908 9722 4936 10066
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 7944 9518 7972 9862
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 16868 9722 16896 10066
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 18432 9518 18460 9862
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 19812 9722 19840 10066
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 26620 9518 26648 9862
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 29564 9722 29592 10066
rect 29552 9716 29604 9722
rect 29552 9658 29604 9664
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8576 9512 8628 9518
rect 12808 9512 12860 9518
rect 8628 9460 8708 9466
rect 8576 9454 8708 9460
rect 12808 9454 12860 9460
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9042 3648 9318
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4724 9178 4752 9454
rect 8588 9438 8708 9454
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 8588 9042 8616 9318
rect 8680 9178 8708 9438
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 7392 8022 7420 8366
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7484 7954 7512 8230
rect 7576 8090 7604 8978
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7760 7954 7788 8230
rect 8036 7954 8064 8774
rect 11164 8634 11192 8978
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11348 8430 11376 9318
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 12820 9178 12848 9454
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 15304 9042 15332 9318
rect 17420 9178 17448 9454
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 22664 9042 22692 9318
rect 23216 9178 23244 9454
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 26528 9042 26556 9318
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 28828 9178 28856 9454
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 29552 9036 29604 9042
rect 29552 8978 29604 8984
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 15120 8430 15148 8774
rect 17880 8634 17908 8978
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8496 7886 8524 8366
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8588 7954 8616 8230
rect 8680 8090 8708 8366
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9048 7954 9076 8230
rect 10704 8090 10732 8366
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 15396 7954 15424 8230
rect 17052 8090 17080 8366
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 18984 7954 19012 8774
rect 19076 8634 19104 8978
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19628 8498 19656 8774
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 21928 8430 21956 8774
rect 22388 8634 22416 8978
rect 24504 8634 24532 8978
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 26712 8430 26740 8774
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 29564 8634 29592 8978
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 24504 8090 24532 8366
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 29104 7954 29132 8230
rect 29288 8090 29316 8366
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 7392 7342 7420 7686
rect 11256 7546 11284 7890
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11348 7426 11376 7686
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 13556 7546 13584 7890
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 11348 7398 11468 7426
rect 11440 7342 11468 7398
rect 15212 7342 15240 7686
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 20364 7546 20392 7890
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 21928 7342 21956 7686
rect 22664 7546 22692 7890
rect 23020 7812 23072 7818
rect 23020 7754 23072 7760
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22756 7342 22784 7686
rect 23032 7342 23060 7754
rect 23492 7478 23520 7890
rect 25976 7546 26004 7890
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 7668 7002 7696 7278
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7760 6866 7788 7142
rect 9968 6866 9996 7142
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 6472 6254 6500 6598
rect 7208 6458 7236 6802
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 10060 6254 10088 6598
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 13464 6458 13492 6802
rect 14108 6798 14136 7278
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6866 15240 7142
rect 17236 7002 17264 7278
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17788 6866 17816 7142
rect 18064 6866 18092 7278
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 6866 18276 7142
rect 19812 7002 19840 7278
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 23492 6934 23520 7142
rect 25792 7002 25820 7278
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 23480 6928 23532 6934
rect 23480 6870 23532 6876
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13648 6254 13676 6598
rect 15948 6458 15976 6802
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 21928 6254 21956 6598
rect 26068 6458 26096 6802
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 5828 5778 5856 6054
rect 8220 5914 8248 6190
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 10244 5778 10272 6054
rect 11164 5914 11192 6190
rect 11716 5914 11744 6190
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11808 5778 11836 6054
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 12636 5778 12664 6054
rect 16684 5914 16712 6190
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 22020 5778 22048 6054
rect 26068 5914 26096 6190
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 6472 5166 6500 5510
rect 9508 5370 9536 5714
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 14292 5166 14320 5510
rect 16408 5370 16436 5714
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 17144 5166 17172 5510
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 19628 5370 19656 5714
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19720 5166 19748 5510
rect 20456 5302 20484 5714
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20732 5234 20760 5510
rect 20824 5370 20852 5714
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 22480 5166 22508 5510
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 7024 4690 7052 4966
rect 9508 4826 9536 5102
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 14936 4690 14964 4966
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 21284 4826 21312 5102
rect 24584 5092 24636 5098
rect 24584 5034 24636 5040
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 24504 4690 24532 4966
rect 24596 4826 24624 5034
rect 24964 4826 24992 5714
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 25608 4690 25636 4966
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 7024 4078 7052 4422
rect 8588 4282 8616 4626
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 11348 4162 11376 4422
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 11900 4282 11928 4626
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11348 4134 11468 4162
rect 11440 4078 11468 4134
rect 12084 4078 12112 4422
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 13832 4026 13860 4626
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15672 4078 15700 4422
rect 17420 4282 17448 4626
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 19628 4078 19656 4422
rect 21836 4282 21864 4626
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 15660 4072 15712 4078
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 6748 3602 6776 3878
rect 8312 3738 8340 4014
rect 13832 3998 13952 4026
rect 15660 4014 15712 4020
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 10244 3602 10272 3878
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 13832 3602 13860 3878
rect 13924 3738 13952 3998
rect 17972 3738 18000 4014
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 20272 3670 20300 3878
rect 24412 3738 24440 4082
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 24504 3602 24532 3878
rect 25148 3738 25176 4014
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25608 3670 25636 3878
rect 25792 3738 25820 4014
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 26160 3602 26188 3878
rect 26896 3738 26924 4014
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 6932 2990 6960 3334
rect 8404 3194 8432 3538
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8680 2990 8708 3334
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 12636 3194 12664 3538
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12912 2990 12940 3334
rect 13004 3194 13032 3538
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13372 2990 13400 3334
rect 18064 3194 18092 3538
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 19720 2990 19748 3334
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 27540 3194 27568 3538
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 7576 2514 7604 2790
rect 11072 2650 11100 2926
rect 11624 2650 11652 2926
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11716 2514 11744 2790
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 13740 2514 13768 2790
rect 13832 2650 13860 2790
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14292 2514 14320 2790
rect 15856 2650 15884 2926
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 18800 2514 18828 2790
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19870 2683 20178 2692
rect 20732 2650 20760 2926
rect 23940 2848 23992 2854
rect 23940 2790 23992 2796
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 23952 2514 23980 2790
rect 26528 2650 26556 2926
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 9048 1902 9076 2246
rect 10428 1970 10456 2246
rect 11072 2106 11100 2450
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11256 2106 11284 2382
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 13556 1902 13584 2246
rect 15580 2106 15608 2450
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 8680 1426 8708 1702
rect 10888 1562 10916 1838
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 13188 1426 13216 1702
rect 16316 1562 16344 1838
rect 18616 1834 18644 2246
rect 19210 2204 19518 2213
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 20640 2106 20668 2450
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 18604 1828 18656 1834
rect 18604 1770 18656 1776
rect 17224 1760 17276 1766
rect 17224 1702 17276 1708
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 17236 1426 17264 1702
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 21100 1494 21128 1906
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 21088 1488 21140 1494
rect 21088 1430 21140 1436
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 13176 1420 13228 1426
rect 13176 1362 13228 1368
rect 16396 1420 16448 1426
rect 16396 1362 16448 1368
rect 17224 1420 17276 1426
rect 17224 1362 17276 1368
rect 18696 1420 18748 1426
rect 18696 1362 18748 1368
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 8956 814 8984 1158
rect 10244 1018 10272 1362
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 10232 1012 10284 1018
rect 10232 954 10284 960
rect 13924 882 13952 1158
rect 16408 1018 16436 1362
rect 17316 1216 17368 1222
rect 17316 1158 17368 1164
rect 16396 1012 16448 1018
rect 16396 954 16448 960
rect 13912 876 13964 882
rect 13912 818 13964 824
rect 17328 814 17356 1158
rect 18708 1018 18736 1362
rect 19892 1216 19944 1222
rect 19892 1158 19944 1164
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 18696 1012 18748 1018
rect 18696 954 18748 960
rect 19904 814 19932 1158
rect 20732 1018 20760 1362
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 20720 1012 20772 1018
rect 20720 954 20772 960
rect 8944 808 8996 814
rect 8944 750 8996 756
rect 17316 808 17368 814
rect 17316 750 17368 756
rect 19892 808 19944 814
rect 19892 750 19944 756
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
<< via2 >>
rect 28630 22072 28686 22128
rect 11794 21936 11850 21992
rect 12254 21936 12310 21992
rect 19706 21936 19762 21992
rect 20350 21936 20406 21992
rect 22650 21936 22706 21992
rect 27526 21936 27582 21992
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 11442 21786 11498 21788
rect 11522 21786 11578 21788
rect 11602 21786 11658 21788
rect 11682 21786 11738 21788
rect 11442 21734 11488 21786
rect 11488 21734 11498 21786
rect 11522 21734 11552 21786
rect 11552 21734 11564 21786
rect 11564 21734 11578 21786
rect 11602 21734 11616 21786
rect 11616 21734 11628 21786
rect 11628 21734 11658 21786
rect 11682 21734 11692 21786
rect 11692 21734 11738 21786
rect 11442 21732 11498 21734
rect 11522 21732 11578 21734
rect 11602 21732 11658 21734
rect 11682 21732 11738 21734
rect 6182 21684 6238 21720
rect 6182 21664 6184 21684
rect 6184 21664 6236 21684
rect 6236 21664 6238 21684
rect 6734 21684 6790 21720
rect 6734 21664 6736 21684
rect 6736 21664 6788 21684
rect 6788 21664 6790 21684
rect 7286 21684 7342 21720
rect 7286 21664 7288 21684
rect 7288 21664 7340 21684
rect 7340 21664 7342 21684
rect 7838 21684 7894 21720
rect 7838 21664 7840 21684
rect 7840 21664 7892 21684
rect 7892 21664 7894 21684
rect 8390 21684 8446 21720
rect 8390 21664 8392 21684
rect 8392 21664 8444 21684
rect 8444 21664 8446 21684
rect 8942 21684 8998 21720
rect 8942 21664 8944 21684
rect 8944 21664 8996 21684
rect 8996 21664 8998 21684
rect 9494 21684 9550 21720
rect 9494 21664 9496 21684
rect 9496 21664 9548 21684
rect 9548 21664 9550 21684
rect 10046 21684 10102 21720
rect 10046 21664 10048 21684
rect 10048 21664 10100 21684
rect 10100 21664 10102 21684
rect 10598 21684 10654 21720
rect 10598 21664 10600 21684
rect 10600 21664 10652 21684
rect 10652 21664 10654 21684
rect 11150 21684 11206 21720
rect 16762 21800 16818 21856
rect 11150 21664 11152 21684
rect 11152 21664 11204 21684
rect 11204 21664 11206 21684
rect 12806 21684 12862 21720
rect 12806 21664 12808 21684
rect 12808 21664 12860 21684
rect 12860 21664 12862 21684
rect 13542 21684 13598 21720
rect 13542 21664 13544 21684
rect 13544 21664 13596 21684
rect 13596 21664 13598 21684
rect 13910 21684 13966 21720
rect 13910 21664 13912 21684
rect 13912 21664 13964 21684
rect 13964 21664 13966 21684
rect 14462 21684 14518 21720
rect 14462 21664 14464 21684
rect 14464 21664 14516 21684
rect 14516 21664 14518 21684
rect 15198 21684 15254 21720
rect 15198 21664 15200 21684
rect 15200 21664 15252 21684
rect 15252 21664 15254 21684
rect 15658 21684 15714 21720
rect 15658 21664 15660 21684
rect 15660 21664 15712 21684
rect 15712 21664 15714 21684
rect 16118 21684 16174 21720
rect 16118 21664 16120 21684
rect 16120 21664 16172 21684
rect 16172 21664 16174 21684
rect 16946 21684 17002 21720
rect 16946 21664 16948 21684
rect 16948 21664 17000 21684
rect 17000 21664 17002 21684
rect 17590 21684 17646 21720
rect 17590 21664 17592 21684
rect 17592 21664 17644 21684
rect 17644 21664 17646 21684
rect 18326 21684 18382 21720
rect 18326 21664 18328 21684
rect 18328 21664 18380 21684
rect 18380 21664 18382 21684
rect 19216 21786 19272 21788
rect 19296 21786 19352 21788
rect 19376 21786 19432 21788
rect 19456 21786 19512 21788
rect 19216 21734 19262 21786
rect 19262 21734 19272 21786
rect 19296 21734 19326 21786
rect 19326 21734 19338 21786
rect 19338 21734 19352 21786
rect 19376 21734 19390 21786
rect 19390 21734 19402 21786
rect 19402 21734 19432 21786
rect 19456 21734 19466 21786
rect 19466 21734 19512 21786
rect 19216 21732 19272 21734
rect 19296 21732 19352 21734
rect 19376 21732 19432 21734
rect 19456 21732 19512 21734
rect 19338 21564 19340 21584
rect 19340 21564 19392 21584
rect 19392 21564 19394 21584
rect 19338 21528 19394 21564
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 12102 21242 12158 21244
rect 12182 21242 12238 21244
rect 12262 21242 12318 21244
rect 12342 21242 12398 21244
rect 12102 21190 12148 21242
rect 12148 21190 12158 21242
rect 12182 21190 12212 21242
rect 12212 21190 12224 21242
rect 12224 21190 12238 21242
rect 12262 21190 12276 21242
rect 12276 21190 12288 21242
rect 12288 21190 12318 21242
rect 12342 21190 12352 21242
rect 12352 21190 12398 21242
rect 12102 21188 12158 21190
rect 12182 21188 12238 21190
rect 12262 21188 12318 21190
rect 12342 21188 12398 21190
rect 20718 21800 20774 21856
rect 22098 21800 22154 21856
rect 21546 21528 21602 21584
rect 19876 21242 19932 21244
rect 19956 21242 20012 21244
rect 20036 21242 20092 21244
rect 20116 21242 20172 21244
rect 19876 21190 19922 21242
rect 19922 21190 19932 21242
rect 19956 21190 19986 21242
rect 19986 21190 19998 21242
rect 19998 21190 20012 21242
rect 20036 21190 20050 21242
rect 20050 21190 20062 21242
rect 20062 21190 20092 21242
rect 20116 21190 20126 21242
rect 20126 21190 20172 21242
rect 19876 21188 19932 21190
rect 19956 21188 20012 21190
rect 20036 21188 20092 21190
rect 20116 21188 20172 21190
rect 22742 21800 22798 21856
rect 24858 21800 24914 21856
rect 23478 21528 23534 21584
rect 24030 21528 24086 21584
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 11442 20698 11498 20700
rect 11522 20698 11578 20700
rect 11602 20698 11658 20700
rect 11682 20698 11738 20700
rect 11442 20646 11488 20698
rect 11488 20646 11498 20698
rect 11522 20646 11552 20698
rect 11552 20646 11564 20698
rect 11564 20646 11578 20698
rect 11602 20646 11616 20698
rect 11616 20646 11628 20698
rect 11628 20646 11658 20698
rect 11682 20646 11692 20698
rect 11692 20646 11738 20698
rect 11442 20644 11498 20646
rect 11522 20644 11578 20646
rect 11602 20644 11658 20646
rect 11682 20644 11738 20646
rect 19216 20698 19272 20700
rect 19296 20698 19352 20700
rect 19376 20698 19432 20700
rect 19456 20698 19512 20700
rect 19216 20646 19262 20698
rect 19262 20646 19272 20698
rect 19296 20646 19326 20698
rect 19326 20646 19338 20698
rect 19338 20646 19352 20698
rect 19376 20646 19390 20698
rect 19390 20646 19402 20698
rect 19402 20646 19432 20698
rect 19456 20646 19466 20698
rect 19466 20646 19512 20698
rect 19216 20644 19272 20646
rect 19296 20644 19352 20646
rect 19376 20644 19432 20646
rect 19456 20644 19512 20646
rect 26990 21786 27046 21788
rect 27070 21786 27126 21788
rect 27150 21786 27206 21788
rect 27230 21786 27286 21788
rect 26990 21734 27036 21786
rect 27036 21734 27046 21786
rect 27070 21734 27100 21786
rect 27100 21734 27112 21786
rect 27112 21734 27126 21786
rect 27150 21734 27164 21786
rect 27164 21734 27176 21786
rect 27176 21734 27206 21786
rect 27230 21734 27240 21786
rect 27240 21734 27286 21786
rect 26990 21732 27046 21734
rect 27070 21732 27126 21734
rect 27150 21732 27206 21734
rect 27230 21732 27286 21734
rect 24950 21528 25006 21584
rect 27250 21528 27306 21584
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 12102 20154 12158 20156
rect 12182 20154 12238 20156
rect 12262 20154 12318 20156
rect 12342 20154 12398 20156
rect 12102 20102 12148 20154
rect 12148 20102 12158 20154
rect 12182 20102 12212 20154
rect 12212 20102 12224 20154
rect 12224 20102 12238 20154
rect 12262 20102 12276 20154
rect 12276 20102 12288 20154
rect 12288 20102 12318 20154
rect 12342 20102 12352 20154
rect 12352 20102 12398 20154
rect 12102 20100 12158 20102
rect 12182 20100 12238 20102
rect 12262 20100 12318 20102
rect 12342 20100 12398 20102
rect 19876 20154 19932 20156
rect 19956 20154 20012 20156
rect 20036 20154 20092 20156
rect 20116 20154 20172 20156
rect 19876 20102 19922 20154
rect 19922 20102 19932 20154
rect 19956 20102 19986 20154
rect 19986 20102 19998 20154
rect 19998 20102 20012 20154
rect 20036 20102 20050 20154
rect 20050 20102 20062 20154
rect 20062 20102 20092 20154
rect 20116 20102 20126 20154
rect 20126 20102 20172 20154
rect 19876 20100 19932 20102
rect 19956 20100 20012 20102
rect 20036 20100 20092 20102
rect 20116 20100 20172 20102
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 11442 19610 11498 19612
rect 11522 19610 11578 19612
rect 11602 19610 11658 19612
rect 11682 19610 11738 19612
rect 11442 19558 11488 19610
rect 11488 19558 11498 19610
rect 11522 19558 11552 19610
rect 11552 19558 11564 19610
rect 11564 19558 11578 19610
rect 11602 19558 11616 19610
rect 11616 19558 11628 19610
rect 11628 19558 11658 19610
rect 11682 19558 11692 19610
rect 11692 19558 11738 19610
rect 11442 19556 11498 19558
rect 11522 19556 11578 19558
rect 11602 19556 11658 19558
rect 11682 19556 11738 19558
rect 19216 19610 19272 19612
rect 19296 19610 19352 19612
rect 19376 19610 19432 19612
rect 19456 19610 19512 19612
rect 19216 19558 19262 19610
rect 19262 19558 19272 19610
rect 19296 19558 19326 19610
rect 19326 19558 19338 19610
rect 19338 19558 19352 19610
rect 19376 19558 19390 19610
rect 19390 19558 19402 19610
rect 19402 19558 19432 19610
rect 19456 19558 19466 19610
rect 19466 19558 19512 19610
rect 19216 19556 19272 19558
rect 19296 19556 19352 19558
rect 19376 19556 19432 19558
rect 19456 19556 19512 19558
rect 27650 21242 27706 21244
rect 27730 21242 27786 21244
rect 27810 21242 27866 21244
rect 27890 21242 27946 21244
rect 27650 21190 27696 21242
rect 27696 21190 27706 21242
rect 27730 21190 27760 21242
rect 27760 21190 27772 21242
rect 27772 21190 27786 21242
rect 27810 21190 27824 21242
rect 27824 21190 27836 21242
rect 27836 21190 27866 21242
rect 27890 21190 27900 21242
rect 27900 21190 27946 21242
rect 27650 21188 27706 21190
rect 27730 21188 27786 21190
rect 27810 21188 27866 21190
rect 27890 21188 27946 21190
rect 29734 21800 29790 21856
rect 28814 21528 28870 21584
rect 26990 20698 27046 20700
rect 27070 20698 27126 20700
rect 27150 20698 27206 20700
rect 27230 20698 27286 20700
rect 26990 20646 27036 20698
rect 27036 20646 27046 20698
rect 27070 20646 27100 20698
rect 27100 20646 27112 20698
rect 27112 20646 27126 20698
rect 27150 20646 27164 20698
rect 27164 20646 27176 20698
rect 27176 20646 27206 20698
rect 27230 20646 27240 20698
rect 27240 20646 27286 20698
rect 26990 20644 27046 20646
rect 27070 20644 27126 20646
rect 27150 20644 27206 20646
rect 27230 20644 27286 20646
rect 26330 19488 26386 19544
rect 26238 19352 26294 19408
rect 27650 20154 27706 20156
rect 27730 20154 27786 20156
rect 27810 20154 27866 20156
rect 27890 20154 27946 20156
rect 27650 20102 27696 20154
rect 27696 20102 27706 20154
rect 27730 20102 27760 20154
rect 27760 20102 27772 20154
rect 27772 20102 27786 20154
rect 27810 20102 27824 20154
rect 27824 20102 27836 20154
rect 27836 20102 27866 20154
rect 27890 20102 27900 20154
rect 27900 20102 27946 20154
rect 27650 20100 27706 20102
rect 27730 20100 27786 20102
rect 27810 20100 27866 20102
rect 27890 20100 27946 20102
rect 26990 19610 27046 19612
rect 27070 19610 27126 19612
rect 27150 19610 27206 19612
rect 27230 19610 27286 19612
rect 26990 19558 27036 19610
rect 27036 19558 27046 19610
rect 27070 19558 27100 19610
rect 27100 19558 27112 19610
rect 27112 19558 27126 19610
rect 27150 19558 27164 19610
rect 27164 19558 27176 19610
rect 27176 19558 27206 19610
rect 27230 19558 27240 19610
rect 27240 19558 27286 19610
rect 26990 19556 27046 19558
rect 27070 19556 27126 19558
rect 27150 19556 27206 19558
rect 27230 19556 27286 19558
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 27654 22068 27660 22132
rect 27724 22130 27730 22132
rect 28625 22130 28691 22133
rect 27724 22128 28691 22130
rect 27724 22072 28630 22128
rect 28686 22072 28691 22128
rect 27724 22070 28691 22072
rect 27724 22068 27730 22070
rect 28625 22067 28691 22070
rect 11646 21932 11652 21996
rect 11716 21994 11722 21996
rect 11789 21994 11855 21997
rect 12249 21996 12315 21997
rect 11716 21992 11855 21994
rect 11716 21936 11794 21992
rect 11850 21936 11855 21992
rect 11716 21934 11855 21936
rect 11716 21932 11722 21934
rect 11789 21931 11855 21934
rect 12198 21932 12204 21996
rect 12268 21994 12315 21996
rect 12268 21992 12360 21994
rect 12310 21936 12360 21992
rect 12268 21934 12360 21936
rect 12268 21932 12315 21934
rect 19374 21932 19380 21996
rect 19444 21994 19450 21996
rect 19701 21994 19767 21997
rect 19444 21992 19767 21994
rect 19444 21936 19706 21992
rect 19762 21936 19767 21992
rect 19444 21934 19767 21936
rect 19444 21932 19450 21934
rect 12249 21931 12315 21932
rect 19701 21931 19767 21934
rect 19926 21932 19932 21996
rect 19996 21994 20002 21996
rect 20345 21994 20411 21997
rect 19996 21992 20411 21994
rect 19996 21936 20350 21992
rect 20406 21936 20411 21992
rect 19996 21934 20411 21936
rect 19996 21932 20002 21934
rect 20345 21931 20411 21934
rect 22134 21932 22140 21996
rect 22204 21994 22210 21996
rect 22645 21994 22711 21997
rect 22204 21992 22711 21994
rect 22204 21936 22650 21992
rect 22706 21936 22711 21992
rect 22204 21934 22711 21936
rect 22204 21932 22210 21934
rect 22645 21931 22711 21934
rect 27102 21932 27108 21996
rect 27172 21994 27178 21996
rect 27521 21994 27587 21997
rect 27172 21992 27587 21994
rect 27172 21936 27526 21992
rect 27582 21936 27587 21992
rect 27172 21934 27587 21936
rect 27172 21932 27178 21934
rect 27521 21931 27587 21934
rect 16757 21858 16823 21861
rect 17166 21858 17172 21860
rect 16757 21856 17172 21858
rect 16757 21800 16762 21856
rect 16818 21800 17172 21856
rect 16757 21798 17172 21800
rect 16757 21795 16823 21798
rect 17166 21796 17172 21798
rect 17236 21796 17242 21860
rect 20478 21796 20484 21860
rect 20548 21858 20554 21860
rect 20713 21858 20779 21861
rect 20548 21856 20779 21858
rect 20548 21800 20718 21856
rect 20774 21800 20779 21856
rect 20548 21798 20779 21800
rect 20548 21796 20554 21798
rect 20713 21795 20779 21798
rect 21582 21796 21588 21860
rect 21652 21858 21658 21860
rect 22093 21858 22159 21861
rect 22737 21860 22803 21861
rect 22686 21858 22692 21860
rect 21652 21856 22159 21858
rect 21652 21800 22098 21856
rect 22154 21800 22159 21856
rect 21652 21798 22159 21800
rect 22646 21798 22692 21858
rect 22756 21856 22803 21860
rect 22798 21800 22803 21856
rect 21652 21796 21658 21798
rect 22093 21795 22159 21798
rect 22686 21796 22692 21798
rect 22756 21796 22803 21800
rect 24342 21796 24348 21860
rect 24412 21858 24418 21860
rect 24853 21858 24919 21861
rect 24412 21856 24919 21858
rect 24412 21800 24858 21856
rect 24914 21800 24919 21856
rect 24412 21798 24919 21800
rect 24412 21796 24418 21798
rect 22737 21795 22803 21796
rect 24853 21795 24919 21798
rect 29310 21796 29316 21860
rect 29380 21858 29386 21860
rect 29729 21858 29795 21861
rect 29380 21856 29795 21858
rect 29380 21800 29734 21856
rect 29790 21800 29795 21856
rect 29380 21798 29795 21800
rect 29380 21796 29386 21798
rect 29729 21795 29795 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 11432 21792 11748 21793
rect 11432 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11748 21792
rect 11432 21727 11748 21728
rect 19206 21792 19522 21793
rect 19206 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19522 21792
rect 19206 21727 19522 21728
rect 26980 21792 27296 21793
rect 26980 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27296 21792
rect 26980 21727 27296 21728
rect 6177 21724 6243 21725
rect 6729 21724 6795 21725
rect 7281 21724 7347 21725
rect 7833 21724 7899 21725
rect 8385 21724 8451 21725
rect 8937 21724 9003 21725
rect 9489 21724 9555 21725
rect 10041 21724 10107 21725
rect 10593 21724 10659 21725
rect 11145 21724 11211 21725
rect 12801 21724 12867 21725
rect 6126 21660 6132 21724
rect 6196 21722 6243 21724
rect 6196 21720 6288 21722
rect 6238 21664 6288 21720
rect 6196 21662 6288 21664
rect 6196 21660 6243 21662
rect 6678 21660 6684 21724
rect 6748 21722 6795 21724
rect 6748 21720 6840 21722
rect 6790 21664 6840 21720
rect 6748 21662 6840 21664
rect 6748 21660 6795 21662
rect 7230 21660 7236 21724
rect 7300 21722 7347 21724
rect 7300 21720 7392 21722
rect 7342 21664 7392 21720
rect 7300 21662 7392 21664
rect 7300 21660 7347 21662
rect 7782 21660 7788 21724
rect 7852 21722 7899 21724
rect 7852 21720 7944 21722
rect 7894 21664 7944 21720
rect 7852 21662 7944 21664
rect 7852 21660 7899 21662
rect 8334 21660 8340 21724
rect 8404 21722 8451 21724
rect 8404 21720 8496 21722
rect 8446 21664 8496 21720
rect 8404 21662 8496 21664
rect 8404 21660 8451 21662
rect 8886 21660 8892 21724
rect 8956 21722 9003 21724
rect 8956 21720 9048 21722
rect 8998 21664 9048 21720
rect 8956 21662 9048 21664
rect 8956 21660 9003 21662
rect 9438 21660 9444 21724
rect 9508 21722 9555 21724
rect 9508 21720 9600 21722
rect 9550 21664 9600 21720
rect 9508 21662 9600 21664
rect 9508 21660 9555 21662
rect 9990 21660 9996 21724
rect 10060 21722 10107 21724
rect 10060 21720 10152 21722
rect 10102 21664 10152 21720
rect 10060 21662 10152 21664
rect 10060 21660 10107 21662
rect 10542 21660 10548 21724
rect 10612 21722 10659 21724
rect 10612 21720 10704 21722
rect 10654 21664 10704 21720
rect 10612 21662 10704 21664
rect 10612 21660 10659 21662
rect 11094 21660 11100 21724
rect 11164 21722 11211 21724
rect 11164 21720 11256 21722
rect 11206 21664 11256 21720
rect 11164 21662 11256 21664
rect 11164 21660 11211 21662
rect 12750 21660 12756 21724
rect 12820 21722 12867 21724
rect 12820 21720 12912 21722
rect 12862 21664 12912 21720
rect 12820 21662 12912 21664
rect 12820 21660 12867 21662
rect 13302 21660 13308 21724
rect 13372 21722 13378 21724
rect 13537 21722 13603 21725
rect 13905 21724 13971 21725
rect 14457 21724 14523 21725
rect 13372 21720 13603 21722
rect 13372 21664 13542 21720
rect 13598 21664 13603 21720
rect 13372 21662 13603 21664
rect 13372 21660 13378 21662
rect 6177 21659 6243 21660
rect 6729 21659 6795 21660
rect 7281 21659 7347 21660
rect 7833 21659 7899 21660
rect 8385 21659 8451 21660
rect 8937 21659 9003 21660
rect 9489 21659 9555 21660
rect 10041 21659 10107 21660
rect 10593 21659 10659 21660
rect 11145 21659 11211 21660
rect 12801 21659 12867 21660
rect 13537 21659 13603 21662
rect 13854 21660 13860 21724
rect 13924 21722 13971 21724
rect 13924 21720 14016 21722
rect 13966 21664 14016 21720
rect 13924 21662 14016 21664
rect 13924 21660 13971 21662
rect 14406 21660 14412 21724
rect 14476 21722 14523 21724
rect 14476 21720 14568 21722
rect 14518 21664 14568 21720
rect 14476 21662 14568 21664
rect 14476 21660 14523 21662
rect 14958 21660 14964 21724
rect 15028 21722 15034 21724
rect 15193 21722 15259 21725
rect 15028 21720 15259 21722
rect 15028 21664 15198 21720
rect 15254 21664 15259 21720
rect 15028 21662 15259 21664
rect 15028 21660 15034 21662
rect 13905 21659 13971 21660
rect 14457 21659 14523 21660
rect 15193 21659 15259 21662
rect 15510 21660 15516 21724
rect 15580 21722 15586 21724
rect 15653 21722 15719 21725
rect 16113 21724 16179 21725
rect 15580 21720 15719 21722
rect 15580 21664 15658 21720
rect 15714 21664 15719 21720
rect 15580 21662 15719 21664
rect 15580 21660 15586 21662
rect 15653 21659 15719 21662
rect 16062 21660 16068 21724
rect 16132 21722 16179 21724
rect 16132 21720 16224 21722
rect 16174 21664 16224 21720
rect 16132 21662 16224 21664
rect 16132 21660 16179 21662
rect 16614 21660 16620 21724
rect 16684 21722 16690 21724
rect 16941 21722 17007 21725
rect 16684 21720 17007 21722
rect 16684 21664 16946 21720
rect 17002 21664 17007 21720
rect 16684 21662 17007 21664
rect 16684 21660 16690 21662
rect 16113 21659 16179 21660
rect 16941 21659 17007 21662
rect 17585 21722 17651 21725
rect 18321 21724 18387 21725
rect 17718 21722 17724 21724
rect 17585 21720 17724 21722
rect 17585 21664 17590 21720
rect 17646 21664 17724 21720
rect 17585 21662 17724 21664
rect 17585 21659 17651 21662
rect 17718 21660 17724 21662
rect 17788 21660 17794 21724
rect 18270 21660 18276 21724
rect 18340 21722 18387 21724
rect 18340 21720 18432 21722
rect 18382 21664 18432 21720
rect 18340 21662 18432 21664
rect 18340 21660 18387 21662
rect 18321 21659 18387 21660
rect 18822 21524 18828 21588
rect 18892 21586 18898 21588
rect 19333 21586 19399 21589
rect 18892 21584 19399 21586
rect 18892 21528 19338 21584
rect 19394 21528 19399 21584
rect 18892 21526 19399 21528
rect 18892 21524 18898 21526
rect 19333 21523 19399 21526
rect 21030 21524 21036 21588
rect 21100 21586 21106 21588
rect 21541 21586 21607 21589
rect 21100 21584 21607 21586
rect 21100 21528 21546 21584
rect 21602 21528 21607 21584
rect 21100 21526 21607 21528
rect 21100 21524 21106 21526
rect 21541 21523 21607 21526
rect 23238 21524 23244 21588
rect 23308 21586 23314 21588
rect 23473 21586 23539 21589
rect 23308 21584 23539 21586
rect 23308 21528 23478 21584
rect 23534 21528 23539 21584
rect 23308 21526 23539 21528
rect 23308 21524 23314 21526
rect 23473 21523 23539 21526
rect 23790 21524 23796 21588
rect 23860 21586 23866 21588
rect 24025 21586 24091 21589
rect 24945 21588 25011 21589
rect 24894 21586 24900 21588
rect 23860 21584 24091 21586
rect 23860 21528 24030 21584
rect 24086 21528 24091 21584
rect 23860 21526 24091 21528
rect 24854 21526 24900 21586
rect 24964 21584 25011 21588
rect 25006 21528 25011 21584
rect 23860 21524 23866 21526
rect 24025 21523 24091 21526
rect 24894 21524 24900 21526
rect 24964 21524 25011 21528
rect 26550 21524 26556 21588
rect 26620 21586 26626 21588
rect 27245 21586 27311 21589
rect 26620 21584 27311 21586
rect 26620 21528 27250 21584
rect 27306 21528 27311 21584
rect 26620 21526 27311 21528
rect 26620 21524 26626 21526
rect 24945 21523 25011 21524
rect 27245 21523 27311 21526
rect 28206 21524 28212 21588
rect 28276 21586 28282 21588
rect 28809 21586 28875 21589
rect 28276 21584 28875 21586
rect 28276 21528 28814 21584
rect 28870 21528 28875 21584
rect 28276 21526 28875 21528
rect 28276 21524 28282 21526
rect 28809 21523 28875 21526
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 12092 21248 12408 21249
rect 12092 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12408 21248
rect 12092 21183 12408 21184
rect 19866 21248 20182 21249
rect 19866 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20182 21248
rect 19866 21183 20182 21184
rect 27640 21248 27956 21249
rect 27640 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27956 21248
rect 27640 21183 27956 21184
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 11432 20704 11748 20705
rect 11432 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11748 20704
rect 11432 20639 11748 20640
rect 19206 20704 19522 20705
rect 19206 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19522 20704
rect 19206 20639 19522 20640
rect 26980 20704 27296 20705
rect 26980 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27296 20704
rect 26980 20639 27296 20640
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 12092 20160 12408 20161
rect 12092 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12408 20160
rect 12092 20095 12408 20096
rect 19866 20160 20182 20161
rect 19866 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20182 20160
rect 19866 20095 20182 20096
rect 27640 20160 27956 20161
rect 27640 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27956 20160
rect 27640 20095 27956 20096
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 11432 19616 11748 19617
rect 11432 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11748 19616
rect 11432 19551 11748 19552
rect 19206 19616 19522 19617
rect 19206 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19522 19616
rect 19206 19551 19522 19552
rect 26980 19616 27296 19617
rect 26980 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27296 19616
rect 26980 19551 27296 19552
rect 25446 19484 25452 19548
rect 25516 19546 25522 19548
rect 26325 19546 26391 19549
rect 25516 19544 26391 19546
rect 25516 19488 26330 19544
rect 26386 19488 26391 19544
rect 25516 19486 26391 19488
rect 25516 19484 25522 19486
rect 26325 19483 26391 19486
rect 25998 19348 26004 19412
rect 26068 19410 26074 19412
rect 26233 19410 26299 19413
rect 26068 19408 26299 19410
rect 26068 19352 26238 19408
rect 26294 19352 26299 19408
rect 26068 19350 26299 19352
rect 26068 19348 26074 19350
rect 26233 19347 26299 19350
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 27660 22068 27724 22132
rect 11652 21932 11716 21996
rect 12204 21992 12268 21996
rect 12204 21936 12254 21992
rect 12254 21936 12268 21992
rect 12204 21932 12268 21936
rect 19380 21932 19444 21996
rect 19932 21932 19996 21996
rect 22140 21932 22204 21996
rect 27108 21932 27172 21996
rect 17172 21796 17236 21860
rect 20484 21796 20548 21860
rect 21588 21796 21652 21860
rect 22692 21856 22756 21860
rect 22692 21800 22742 21856
rect 22742 21800 22756 21856
rect 22692 21796 22756 21800
rect 24348 21796 24412 21860
rect 29316 21796 29380 21860
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 11438 21788 11502 21792
rect 11438 21732 11442 21788
rect 11442 21732 11498 21788
rect 11498 21732 11502 21788
rect 11438 21728 11502 21732
rect 11518 21788 11582 21792
rect 11518 21732 11522 21788
rect 11522 21732 11578 21788
rect 11578 21732 11582 21788
rect 11518 21728 11582 21732
rect 11598 21788 11662 21792
rect 11598 21732 11602 21788
rect 11602 21732 11658 21788
rect 11658 21732 11662 21788
rect 11598 21728 11662 21732
rect 11678 21788 11742 21792
rect 11678 21732 11682 21788
rect 11682 21732 11738 21788
rect 11738 21732 11742 21788
rect 11678 21728 11742 21732
rect 19212 21788 19276 21792
rect 19212 21732 19216 21788
rect 19216 21732 19272 21788
rect 19272 21732 19276 21788
rect 19212 21728 19276 21732
rect 19292 21788 19356 21792
rect 19292 21732 19296 21788
rect 19296 21732 19352 21788
rect 19352 21732 19356 21788
rect 19292 21728 19356 21732
rect 19372 21788 19436 21792
rect 19372 21732 19376 21788
rect 19376 21732 19432 21788
rect 19432 21732 19436 21788
rect 19372 21728 19436 21732
rect 19452 21788 19516 21792
rect 19452 21732 19456 21788
rect 19456 21732 19512 21788
rect 19512 21732 19516 21788
rect 19452 21728 19516 21732
rect 26986 21788 27050 21792
rect 26986 21732 26990 21788
rect 26990 21732 27046 21788
rect 27046 21732 27050 21788
rect 26986 21728 27050 21732
rect 27066 21788 27130 21792
rect 27066 21732 27070 21788
rect 27070 21732 27126 21788
rect 27126 21732 27130 21788
rect 27066 21728 27130 21732
rect 27146 21788 27210 21792
rect 27146 21732 27150 21788
rect 27150 21732 27206 21788
rect 27206 21732 27210 21788
rect 27146 21728 27210 21732
rect 27226 21788 27290 21792
rect 27226 21732 27230 21788
rect 27230 21732 27286 21788
rect 27286 21732 27290 21788
rect 27226 21728 27290 21732
rect 6132 21720 6196 21724
rect 6132 21664 6182 21720
rect 6182 21664 6196 21720
rect 6132 21660 6196 21664
rect 6684 21720 6748 21724
rect 6684 21664 6734 21720
rect 6734 21664 6748 21720
rect 6684 21660 6748 21664
rect 7236 21720 7300 21724
rect 7236 21664 7286 21720
rect 7286 21664 7300 21720
rect 7236 21660 7300 21664
rect 7788 21720 7852 21724
rect 7788 21664 7838 21720
rect 7838 21664 7852 21720
rect 7788 21660 7852 21664
rect 8340 21720 8404 21724
rect 8340 21664 8390 21720
rect 8390 21664 8404 21720
rect 8340 21660 8404 21664
rect 8892 21720 8956 21724
rect 8892 21664 8942 21720
rect 8942 21664 8956 21720
rect 8892 21660 8956 21664
rect 9444 21720 9508 21724
rect 9444 21664 9494 21720
rect 9494 21664 9508 21720
rect 9444 21660 9508 21664
rect 9996 21720 10060 21724
rect 9996 21664 10046 21720
rect 10046 21664 10060 21720
rect 9996 21660 10060 21664
rect 10548 21720 10612 21724
rect 10548 21664 10598 21720
rect 10598 21664 10612 21720
rect 10548 21660 10612 21664
rect 11100 21720 11164 21724
rect 11100 21664 11150 21720
rect 11150 21664 11164 21720
rect 11100 21660 11164 21664
rect 12756 21720 12820 21724
rect 12756 21664 12806 21720
rect 12806 21664 12820 21720
rect 12756 21660 12820 21664
rect 13308 21660 13372 21724
rect 13860 21720 13924 21724
rect 13860 21664 13910 21720
rect 13910 21664 13924 21720
rect 13860 21660 13924 21664
rect 14412 21720 14476 21724
rect 14412 21664 14462 21720
rect 14462 21664 14476 21720
rect 14412 21660 14476 21664
rect 14964 21660 15028 21724
rect 15516 21660 15580 21724
rect 16068 21720 16132 21724
rect 16068 21664 16118 21720
rect 16118 21664 16132 21720
rect 16068 21660 16132 21664
rect 16620 21660 16684 21724
rect 17724 21660 17788 21724
rect 18276 21720 18340 21724
rect 18276 21664 18326 21720
rect 18326 21664 18340 21720
rect 18276 21660 18340 21664
rect 18828 21524 18892 21588
rect 21036 21524 21100 21588
rect 23244 21524 23308 21588
rect 23796 21524 23860 21588
rect 24900 21584 24964 21588
rect 24900 21528 24950 21584
rect 24950 21528 24964 21584
rect 24900 21524 24964 21528
rect 26556 21524 26620 21588
rect 28212 21524 28276 21588
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 12098 21244 12162 21248
rect 12098 21188 12102 21244
rect 12102 21188 12158 21244
rect 12158 21188 12162 21244
rect 12098 21184 12162 21188
rect 12178 21244 12242 21248
rect 12178 21188 12182 21244
rect 12182 21188 12238 21244
rect 12238 21188 12242 21244
rect 12178 21184 12242 21188
rect 12258 21244 12322 21248
rect 12258 21188 12262 21244
rect 12262 21188 12318 21244
rect 12318 21188 12322 21244
rect 12258 21184 12322 21188
rect 12338 21244 12402 21248
rect 12338 21188 12342 21244
rect 12342 21188 12398 21244
rect 12398 21188 12402 21244
rect 12338 21184 12402 21188
rect 19872 21244 19936 21248
rect 19872 21188 19876 21244
rect 19876 21188 19932 21244
rect 19932 21188 19936 21244
rect 19872 21184 19936 21188
rect 19952 21244 20016 21248
rect 19952 21188 19956 21244
rect 19956 21188 20012 21244
rect 20012 21188 20016 21244
rect 19952 21184 20016 21188
rect 20032 21244 20096 21248
rect 20032 21188 20036 21244
rect 20036 21188 20092 21244
rect 20092 21188 20096 21244
rect 20032 21184 20096 21188
rect 20112 21244 20176 21248
rect 20112 21188 20116 21244
rect 20116 21188 20172 21244
rect 20172 21188 20176 21244
rect 20112 21184 20176 21188
rect 27646 21244 27710 21248
rect 27646 21188 27650 21244
rect 27650 21188 27706 21244
rect 27706 21188 27710 21244
rect 27646 21184 27710 21188
rect 27726 21244 27790 21248
rect 27726 21188 27730 21244
rect 27730 21188 27786 21244
rect 27786 21188 27790 21244
rect 27726 21184 27790 21188
rect 27806 21244 27870 21248
rect 27806 21188 27810 21244
rect 27810 21188 27866 21244
rect 27866 21188 27870 21244
rect 27806 21184 27870 21188
rect 27886 21244 27950 21248
rect 27886 21188 27890 21244
rect 27890 21188 27946 21244
rect 27946 21188 27950 21244
rect 27886 21184 27950 21188
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 11438 20700 11502 20704
rect 11438 20644 11442 20700
rect 11442 20644 11498 20700
rect 11498 20644 11502 20700
rect 11438 20640 11502 20644
rect 11518 20700 11582 20704
rect 11518 20644 11522 20700
rect 11522 20644 11578 20700
rect 11578 20644 11582 20700
rect 11518 20640 11582 20644
rect 11598 20700 11662 20704
rect 11598 20644 11602 20700
rect 11602 20644 11658 20700
rect 11658 20644 11662 20700
rect 11598 20640 11662 20644
rect 11678 20700 11742 20704
rect 11678 20644 11682 20700
rect 11682 20644 11738 20700
rect 11738 20644 11742 20700
rect 11678 20640 11742 20644
rect 19212 20700 19276 20704
rect 19212 20644 19216 20700
rect 19216 20644 19272 20700
rect 19272 20644 19276 20700
rect 19212 20640 19276 20644
rect 19292 20700 19356 20704
rect 19292 20644 19296 20700
rect 19296 20644 19352 20700
rect 19352 20644 19356 20700
rect 19292 20640 19356 20644
rect 19372 20700 19436 20704
rect 19372 20644 19376 20700
rect 19376 20644 19432 20700
rect 19432 20644 19436 20700
rect 19372 20640 19436 20644
rect 19452 20700 19516 20704
rect 19452 20644 19456 20700
rect 19456 20644 19512 20700
rect 19512 20644 19516 20700
rect 19452 20640 19516 20644
rect 26986 20700 27050 20704
rect 26986 20644 26990 20700
rect 26990 20644 27046 20700
rect 27046 20644 27050 20700
rect 26986 20640 27050 20644
rect 27066 20700 27130 20704
rect 27066 20644 27070 20700
rect 27070 20644 27126 20700
rect 27126 20644 27130 20700
rect 27066 20640 27130 20644
rect 27146 20700 27210 20704
rect 27146 20644 27150 20700
rect 27150 20644 27206 20700
rect 27206 20644 27210 20700
rect 27146 20640 27210 20644
rect 27226 20700 27290 20704
rect 27226 20644 27230 20700
rect 27230 20644 27286 20700
rect 27286 20644 27290 20700
rect 27226 20640 27290 20644
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 12098 20156 12162 20160
rect 12098 20100 12102 20156
rect 12102 20100 12158 20156
rect 12158 20100 12162 20156
rect 12098 20096 12162 20100
rect 12178 20156 12242 20160
rect 12178 20100 12182 20156
rect 12182 20100 12238 20156
rect 12238 20100 12242 20156
rect 12178 20096 12242 20100
rect 12258 20156 12322 20160
rect 12258 20100 12262 20156
rect 12262 20100 12318 20156
rect 12318 20100 12322 20156
rect 12258 20096 12322 20100
rect 12338 20156 12402 20160
rect 12338 20100 12342 20156
rect 12342 20100 12398 20156
rect 12398 20100 12402 20156
rect 12338 20096 12402 20100
rect 19872 20156 19936 20160
rect 19872 20100 19876 20156
rect 19876 20100 19932 20156
rect 19932 20100 19936 20156
rect 19872 20096 19936 20100
rect 19952 20156 20016 20160
rect 19952 20100 19956 20156
rect 19956 20100 20012 20156
rect 20012 20100 20016 20156
rect 19952 20096 20016 20100
rect 20032 20156 20096 20160
rect 20032 20100 20036 20156
rect 20036 20100 20092 20156
rect 20092 20100 20096 20156
rect 20032 20096 20096 20100
rect 20112 20156 20176 20160
rect 20112 20100 20116 20156
rect 20116 20100 20172 20156
rect 20172 20100 20176 20156
rect 20112 20096 20176 20100
rect 27646 20156 27710 20160
rect 27646 20100 27650 20156
rect 27650 20100 27706 20156
rect 27706 20100 27710 20156
rect 27646 20096 27710 20100
rect 27726 20156 27790 20160
rect 27726 20100 27730 20156
rect 27730 20100 27786 20156
rect 27786 20100 27790 20156
rect 27726 20096 27790 20100
rect 27806 20156 27870 20160
rect 27806 20100 27810 20156
rect 27810 20100 27866 20156
rect 27866 20100 27870 20156
rect 27806 20096 27870 20100
rect 27886 20156 27950 20160
rect 27886 20100 27890 20156
rect 27890 20100 27946 20156
rect 27946 20100 27950 20156
rect 27886 20096 27950 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 11438 19612 11502 19616
rect 11438 19556 11442 19612
rect 11442 19556 11498 19612
rect 11498 19556 11502 19612
rect 11438 19552 11502 19556
rect 11518 19612 11582 19616
rect 11518 19556 11522 19612
rect 11522 19556 11578 19612
rect 11578 19556 11582 19612
rect 11518 19552 11582 19556
rect 11598 19612 11662 19616
rect 11598 19556 11602 19612
rect 11602 19556 11658 19612
rect 11658 19556 11662 19612
rect 11598 19552 11662 19556
rect 11678 19612 11742 19616
rect 11678 19556 11682 19612
rect 11682 19556 11738 19612
rect 11738 19556 11742 19612
rect 11678 19552 11742 19556
rect 19212 19612 19276 19616
rect 19212 19556 19216 19612
rect 19216 19556 19272 19612
rect 19272 19556 19276 19612
rect 19212 19552 19276 19556
rect 19292 19612 19356 19616
rect 19292 19556 19296 19612
rect 19296 19556 19352 19612
rect 19352 19556 19356 19612
rect 19292 19552 19356 19556
rect 19372 19612 19436 19616
rect 19372 19556 19376 19612
rect 19376 19556 19432 19612
rect 19432 19556 19436 19612
rect 19372 19552 19436 19556
rect 19452 19612 19516 19616
rect 19452 19556 19456 19612
rect 19456 19556 19512 19612
rect 19512 19556 19516 19612
rect 19452 19552 19516 19556
rect 26986 19612 27050 19616
rect 26986 19556 26990 19612
rect 26990 19556 27046 19612
rect 27046 19556 27050 19612
rect 26986 19552 27050 19556
rect 27066 19612 27130 19616
rect 27066 19556 27070 19612
rect 27070 19556 27126 19612
rect 27126 19556 27130 19612
rect 27066 19552 27130 19556
rect 27146 19612 27210 19616
rect 27146 19556 27150 19612
rect 27150 19556 27206 19612
rect 27206 19556 27210 19612
rect 27146 19552 27210 19556
rect 27226 19612 27290 19616
rect 27226 19556 27230 19612
rect 27230 19556 27286 19612
rect 27286 19556 27290 19612
rect 27226 19552 27290 19556
rect 25452 19484 25516 19548
rect 26004 19348 26068 19412
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 21792 3976 21808
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 21248 4636 21808
rect 6134 21725 6194 22304
rect 6686 21725 6746 22304
rect 7238 21725 7298 22304
rect 7790 21725 7850 22304
rect 8342 21725 8402 22304
rect 8894 21725 8954 22304
rect 9446 21725 9506 22304
rect 9998 21725 10058 22304
rect 10550 21725 10610 22304
rect 11102 21725 11162 22304
rect 11654 21997 11714 22304
rect 12206 21997 12266 22304
rect 11651 21996 11717 21997
rect 11651 21932 11652 21996
rect 11716 21932 11717 21996
rect 11651 21931 11717 21932
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 11430 21792 11750 21808
rect 11430 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11750 21792
rect 6131 21724 6197 21725
rect 6131 21660 6132 21724
rect 6196 21660 6197 21724
rect 6131 21659 6197 21660
rect 6683 21724 6749 21725
rect 6683 21660 6684 21724
rect 6748 21660 6749 21724
rect 6683 21659 6749 21660
rect 7235 21724 7301 21725
rect 7235 21660 7236 21724
rect 7300 21660 7301 21724
rect 7235 21659 7301 21660
rect 7787 21724 7853 21725
rect 7787 21660 7788 21724
rect 7852 21660 7853 21724
rect 7787 21659 7853 21660
rect 8339 21724 8405 21725
rect 8339 21660 8340 21724
rect 8404 21660 8405 21724
rect 8339 21659 8405 21660
rect 8891 21724 8957 21725
rect 8891 21660 8892 21724
rect 8956 21660 8957 21724
rect 8891 21659 8957 21660
rect 9443 21724 9509 21725
rect 9443 21660 9444 21724
rect 9508 21660 9509 21724
rect 9443 21659 9509 21660
rect 9995 21724 10061 21725
rect 9995 21660 9996 21724
rect 10060 21660 10061 21724
rect 9995 21659 10061 21660
rect 10547 21724 10613 21725
rect 10547 21660 10548 21724
rect 10612 21660 10613 21724
rect 10547 21659 10613 21660
rect 11099 21724 11165 21725
rect 11099 21660 11100 21724
rect 11164 21660 11165 21724
rect 11099 21659 11165 21660
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 20704 11750 21728
rect 11430 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11750 20704
rect 11430 19616 11750 20640
rect 11430 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11750 19616
rect 11430 18528 11750 19552
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 11430 17440 11750 18464
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11430 16352 11750 17376
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11430 15264 11750 16288
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11430 8736 11750 9760
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 21248 12410 21808
rect 12758 21725 12818 22304
rect 13310 21725 13370 22304
rect 13862 21725 13922 22304
rect 14414 21725 14474 22304
rect 14966 21725 15026 22304
rect 15518 21725 15578 22304
rect 16070 21725 16130 22304
rect 16622 21725 16682 22304
rect 17174 21861 17234 22304
rect 17171 21860 17237 21861
rect 17171 21796 17172 21860
rect 17236 21796 17237 21860
rect 17171 21795 17237 21796
rect 17726 21725 17786 22304
rect 18278 21725 18338 22304
rect 12755 21724 12821 21725
rect 12755 21660 12756 21724
rect 12820 21660 12821 21724
rect 12755 21659 12821 21660
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 13859 21724 13925 21725
rect 13859 21660 13860 21724
rect 13924 21660 13925 21724
rect 13859 21659 13925 21660
rect 14411 21724 14477 21725
rect 14411 21660 14412 21724
rect 14476 21660 14477 21724
rect 14411 21659 14477 21660
rect 14963 21724 15029 21725
rect 14963 21660 14964 21724
rect 15028 21660 15029 21724
rect 14963 21659 15029 21660
rect 15515 21724 15581 21725
rect 15515 21660 15516 21724
rect 15580 21660 15581 21724
rect 15515 21659 15581 21660
rect 16067 21724 16133 21725
rect 16067 21660 16068 21724
rect 16132 21660 16133 21724
rect 16067 21659 16133 21660
rect 16619 21724 16685 21725
rect 16619 21660 16620 21724
rect 16684 21660 16685 21724
rect 16619 21659 16685 21660
rect 17723 21724 17789 21725
rect 17723 21660 17724 21724
rect 17788 21660 17789 21724
rect 17723 21659 17789 21660
rect 18275 21724 18341 21725
rect 18275 21660 18276 21724
rect 18340 21660 18341 21724
rect 18275 21659 18341 21660
rect 18830 21589 18890 22304
rect 19382 21997 19442 22304
rect 19934 21997 19994 22304
rect 19379 21996 19445 21997
rect 19379 21932 19380 21996
rect 19444 21932 19445 21996
rect 19379 21931 19445 21932
rect 19931 21996 19997 21997
rect 19931 21932 19932 21996
rect 19996 21932 19997 21996
rect 19931 21931 19997 21932
rect 20486 21861 20546 22304
rect 20483 21860 20549 21861
rect 19204 21792 19524 21808
rect 19204 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19524 21792
rect 18827 21588 18893 21589
rect 18827 21524 18828 21588
rect 18892 21524 18893 21588
rect 18827 21523 18893 21524
rect 12090 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12410 21248
rect 12090 20160 12410 21184
rect 12090 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12410 20160
rect 12090 19072 12410 20096
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 12090 17984 12410 19008
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 12090 16896 12410 17920
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 12090 15808 12410 16832
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 12090 14720 12410 15744
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 20704 19524 21728
rect 19204 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19524 20704
rect 19204 19616 19524 20640
rect 19204 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19524 19616
rect 19204 18528 19524 19552
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 21248 20184 21808
rect 20483 21796 20484 21860
rect 20548 21796 20549 21860
rect 20483 21795 20549 21796
rect 21038 21589 21098 22304
rect 21590 21861 21650 22304
rect 22142 21997 22202 22304
rect 22139 21996 22205 21997
rect 22139 21932 22140 21996
rect 22204 21932 22205 21996
rect 22139 21931 22205 21932
rect 22694 21861 22754 22304
rect 21587 21860 21653 21861
rect 21587 21796 21588 21860
rect 21652 21796 21653 21860
rect 21587 21795 21653 21796
rect 22691 21860 22757 21861
rect 22691 21796 22692 21860
rect 22756 21796 22757 21860
rect 22691 21795 22757 21796
rect 23246 21589 23306 22304
rect 23798 21589 23858 22304
rect 24350 21861 24410 22304
rect 24347 21860 24413 21861
rect 24347 21796 24348 21860
rect 24412 21796 24413 21860
rect 24347 21795 24413 21796
rect 24902 21589 24962 22304
rect 21035 21588 21101 21589
rect 21035 21524 21036 21588
rect 21100 21524 21101 21588
rect 21035 21523 21101 21524
rect 23243 21588 23309 21589
rect 23243 21524 23244 21588
rect 23308 21524 23309 21588
rect 23243 21523 23309 21524
rect 23795 21588 23861 21589
rect 23795 21524 23796 21588
rect 23860 21524 23861 21588
rect 23795 21523 23861 21524
rect 24899 21588 24965 21589
rect 24899 21524 24900 21588
rect 24964 21524 24965 21588
rect 24899 21523 24965 21524
rect 19864 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20184 21248
rect 19864 20160 20184 21184
rect 19864 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20184 20160
rect 19864 19072 20184 20096
rect 25454 19549 25514 22304
rect 25451 19548 25517 19549
rect 25451 19484 25452 19548
rect 25516 19484 25517 19548
rect 25451 19483 25517 19484
rect 26006 19413 26066 22304
rect 26558 21589 26618 22304
rect 27110 21997 27170 22304
rect 27662 22133 27722 22304
rect 27659 22132 27725 22133
rect 27659 22068 27660 22132
rect 27724 22068 27725 22132
rect 27659 22067 27725 22068
rect 27107 21996 27173 21997
rect 27107 21932 27108 21996
rect 27172 21932 27173 21996
rect 27107 21931 27173 21932
rect 26978 21792 27298 21808
rect 26978 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27298 21792
rect 26555 21588 26621 21589
rect 26555 21524 26556 21588
rect 26620 21524 26621 21588
rect 26555 21523 26621 21524
rect 26978 20704 27298 21728
rect 26978 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27298 20704
rect 26978 19616 27298 20640
rect 26978 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27298 19616
rect 26003 19412 26069 19413
rect 26003 19348 26004 19412
rect 26068 19348 26069 19412
rect 26003 19347 26069 19348
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19864 10368 20184 11392
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 18528 27298 19552
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 26978 15264 27298 16288
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26978 7648 27298 8672
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 21248 27958 21808
rect 28214 21589 28274 22304
rect 28766 22104 28826 22304
rect 29318 21861 29378 22304
rect 29315 21860 29381 21861
rect 29315 21796 29316 21860
rect 29380 21796 29381 21860
rect 29315 21795 29381 21796
rect 28211 21588 28277 21589
rect 28211 21524 28212 21588
rect 28276 21524 28277 21588
rect 28211 21523 28277 21524
rect 27638 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27958 21248
rect 27638 20160 27958 21184
rect 27638 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27958 20160
rect 27638 19072 27958 20096
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27638 14720 27958 15744
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27638 7104 27958 8128
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__and4_1  _05_
timestamp 1
transform -1 0 26036 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _06_
timestamp 1
transform 1 0 23092 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _07_
timestamp 1
transform -1 0 22172 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _08_
timestamp 1
transform 1 0 23828 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _09_
timestamp 1
transform 1 0 24472 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _10_
timestamp 1
transform -1 0 27048 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1
transform -1 0 19688 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1
transform -1 0 18584 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1
transform 1 0 17388 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1
transform 1 0 16560 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1
transform -1 0 15640 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_104
timestamp 1
transform 1 0 10120 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1
transform 1 0 13524 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_161
timestamp 1
transform 1 0 15364 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1
transform 1 0 16100 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_177
timestamp 1
transform 1 0 16836 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_200
timestamp 1
transform 1 0 18952 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_211
timestamp 1
transform 1 0 19964 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 1
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_81
timestamp 1
transform 1 0 8004 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1
transform 1 0 8556 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_100
timestamp 1
transform 1 0 9752 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1
transform 1 0 10948 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_123
timestamp 1636968456
transform 1 0 11868 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_135
timestamp 1
transform 1 0 12972 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_161
timestamp 1
transform 1 0 15364 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1
transform 1 0 15824 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_175
timestamp 1
transform 1 0 16652 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_188
timestamp 1
transform 1 0 17848 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_196
timestamp 1
transform 1 0 18584 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_212
timestamp 1
transform 1 0 20056 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_216
timestamp 1
transform 1 0 20424 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_231
timestamp 1636968456
transform 1 0 21804 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_243
timestamp 1636968456
transform 1 0 22908 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_255
timestamp 1636968456
transform 1 0 24012 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_267
timestamp 1636968456
transform 1 0 25116 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1
transform 1 0 30820 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1
transform 1 0 8372 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_99
timestamp 1
transform 1 0 9660 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_107
timestamp 1
transform 1 0 10396 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_125
timestamp 1
transform 1 0 12052 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_147
timestamp 1636968456
transform 1 0 14076 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_159
timestamp 1
transform 1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_174
timestamp 1
transform 1 0 16560 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_206
timestamp 1
transform 1 0 19504 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_214
timestamp 1
transform 1 0 20240 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_229
timestamp 1636968456
transform 1 0 21620 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1
transform 1 0 22724 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1
transform 1 0 23460 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_88
timestamp 1
transform 1 0 8648 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_98
timestamp 1
transform 1 0 9568 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_124
timestamp 1636968456
transform 1 0 11960 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_136
timestamp 1
transform 1 0 13064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_146
timestamp 1
transform 1 0 13984 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_153
timestamp 1
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_161
timestamp 1
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_175
timestamp 1636968456
transform 1 0 16652 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_187
timestamp 1
transform 1 0 17756 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_207
timestamp 1
transform 1 0 19596 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_228
timestamp 1636968456
transform 1 0 21528 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_240
timestamp 1636968456
transform 1 0 22632 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_290
timestamp 1636968456
transform 1 0 27232 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_302
timestamp 1636968456
transform 1 0 28336 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_314
timestamp 1636968456
transform 1 0 29440 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_326
timestamp 1
transform 1 0 30544 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_334
timestamp 1
transform 1 0 31280 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1
transform 1 0 5428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_61
timestamp 1
transform 1 0 6164 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_73
timestamp 1
transform 1 0 7268 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_91
timestamp 1636968456
transform 1 0 8924 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_103
timestamp 1
transform 1 0 10028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_111
timestamp 1
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_133
timestamp 1
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_158
timestamp 1
transform 1 0 15088 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_188
timestamp 1
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_192
timestamp 1
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_211
timestamp 1
transform 1 0 19964 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_262
timestamp 1636968456
transform 1 0 24656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_274
timestamp 1
transform 1 0 25760 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_292
timestamp 1636968456
transform 1 0 27416 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_304
timestamp 1
transform 1 0 28520 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636968456
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636968456
transform 1 0 30084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 1
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_79
timestamp 1
transform 1 0 7820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_104
timestamp 1
transform 1 0 10120 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_125
timestamp 1
transform 1 0 12052 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_131
timestamp 1
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_135
timestamp 1
transform 1 0 12972 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_141
timestamp 1
transform 1 0 13524 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_147
timestamp 1636968456
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_159
timestamp 1
transform 1 0 15180 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636968456
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_201
timestamp 1
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_218
timestamp 1
transform 1 0 20608 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_249
timestamp 1
transform 1 0 23460 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_257
timestamp 1
transform 1 0 24196 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_264
timestamp 1
transform 1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_270
timestamp 1
transform 1 0 25392 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_296
timestamp 1636968456
transform 1 0 27784 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_308
timestamp 1636968456
transform 1 0 28888 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_320
timestamp 1636968456
transform 1 0 29992 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_332
timestamp 1
transform 1 0 31096 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_77
timestamp 1
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_96
timestamp 1
transform 1 0 9384 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_102
timestamp 1
transform 1 0 9936 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_121
timestamp 1
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_128
timestamp 1636968456
transform 1 0 12328 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_173
timestamp 1
transform 1 0 16468 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_181
timestamp 1
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_197
timestamp 1
transform 1 0 18676 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_217
timestamp 1
transform 1 0 20516 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636968456
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636968456
transform 1 0 30084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1
transform 1 0 5796 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1
transform 1 0 6532 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_80
timestamp 1
transform 1 0 7912 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_86
timestamp 1
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_99
timestamp 1636968456
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 1
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_137
timestamp 1
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_148
timestamp 1
transform 1 0 14168 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_162
timestamp 1
transform 1 0 15456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_172
timestamp 1
transform 1 0 16376 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_180
timestamp 1
transform 1 0 17112 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_213
timestamp 1
transform 1 0 20148 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_234
timestamp 1636968456
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_246
timestamp 1636968456
transform 1 0 23184 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_261
timestamp 1
transform 1 0 24564 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_267
timestamp 1636968456
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636968456
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636968456
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1
transform 1 0 30820 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636968456
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636968456
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_53
timestamp 1
transform 1 0 5428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_61
timestamp 1
transform 1 0 6164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1
transform 1 0 7544 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1
transform 1 0 8372 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_100
timestamp 1636968456
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_112
timestamp 1636968456
transform 1 0 10856 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_124
timestamp 1636968456
transform 1 0 11960 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 1
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp 1
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_161
timestamp 1
transform 1 0 15364 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_165
timestamp 1
transform 1 0 15732 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_181
timestamp 1636968456
transform 1 0 17204 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1
transform 1 0 18308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_200
timestamp 1
transform 1 0 18952 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_208
timestamp 1
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_212
timestamp 1
transform 1 0 20056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_228
timestamp 1
transform 1 0 21528 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_274
timestamp 1636968456
transform 1 0 25760 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_286
timestamp 1636968456
transform 1 0 26864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_298
timestamp 1
transform 1 0 27968 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1
transform 1 0 28704 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1636968456
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1636968456
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_333
timestamp 1
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636968456
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636968456
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_51
timestamp 1
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_68
timestamp 1636968456
transform 1 0 6808 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_80
timestamp 1
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_125
timestamp 1
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_147
timestamp 1
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_154
timestamp 1
transform 1 0 14720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_162
timestamp 1
transform 1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_175
timestamp 1
transform 1 0 16652 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_179
timestamp 1
transform 1 0 17020 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_225
timestamp 1
transform 1 0 21252 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_243
timestamp 1636968456
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_255
timestamp 1
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_263
timestamp 1
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp 1
transform 1 0 26036 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636968456
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1636968456
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636968456
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636968456
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_53
timestamp 1
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_68
timestamp 1
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_88
timestamp 1636968456
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_100
timestamp 1
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_109
timestamp 1
transform 1 0 10580 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_131
timestamp 1
transform 1 0 12604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1
transform 1 0 13524 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_145
timestamp 1636968456
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_157
timestamp 1
transform 1 0 14996 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 1
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_178
timestamp 1636968456
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1
transform 1 0 18032 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_221
timestamp 1
transform 1 0 20884 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_242
timestamp 1
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1
transform 1 0 23552 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636968456
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_265
timestamp 1
transform 1 0 24932 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_280
timestamp 1636968456
transform 1 0 26312 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_292
timestamp 1636968456
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 1
transform 1 0 28520 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1636968456
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1636968456
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_333
timestamp 1
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636968456
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1
transform 1 0 5796 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_73
timestamp 1
transform 1 0 7268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_77
timestamp 1
transform 1 0 7636 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636968456
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_93
timestamp 1
transform 1 0 9108 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636968456
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636968456
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_137
timestamp 1
transform 1 0 13156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_156
timestamp 1
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_163
timestamp 1
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_185
timestamp 1
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_190
timestamp 1
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_195
timestamp 1
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_214
timestamp 1
transform 1 0 20240 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1
transform 1 0 20976 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_225
timestamp 1
transform 1 0 21252 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1636968456
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_261
timestamp 1
transform 1 0 24564 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_267
timestamp 1
transform 1 0 25116 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636968456
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636968456
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636968456
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1636968456
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1
transform 1 0 30820 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636968456
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_65
timestamp 1
transform 1 0 6532 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_106
timestamp 1
transform 1 0 10304 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_114
timestamp 1
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636968456
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_150
timestamp 1
transform 1 0 14352 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_158
timestamp 1
transform 1 0 15088 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_168
timestamp 1636968456
transform 1 0 16008 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_189
timestamp 1
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_197
timestamp 1
transform 1 0 18676 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_205
timestamp 1
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_219
timestamp 1
transform 1 0 20700 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_227
timestamp 1
transform 1 0 21436 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_233
timestamp 1
transform 1 0 21988 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_265
timestamp 1
transform 1 0 24932 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1636968456
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1636968456
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1636968456
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636968456
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636968456
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636968456
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_69
timestamp 1
transform 1 0 6900 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_90
timestamp 1
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_95
timestamp 1636968456
transform 1 0 9292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_107
timestamp 1
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_145
timestamp 1
transform 1 0 13892 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_153
timestamp 1
transform 1 0 14628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_172
timestamp 1
transform 1 0 16376 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_201
timestamp 1636968456
transform 1 0 19044 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1
transform 1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_252
timestamp 1
transform 1 0 23736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_311
timestamp 1636968456
transform 1 0 29164 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_323
timestamp 1636968456
transform 1 0 30268 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636968456
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636968456
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636968456
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_65
timestamp 1
transform 1 0 6532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_71
timestamp 1
transform 1 0 7084 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_113
timestamp 1
transform 1 0 10948 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_117
timestamp 1
transform 1 0 11316 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1636968456
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636968456
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_170
timestamp 1
transform 1 0 16192 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_176
timestamp 1
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_197
timestamp 1
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_211
timestamp 1636968456
transform 1 0 19964 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_223
timestamp 1
transform 1 0 21068 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_229
timestamp 1
transform 1 0 21620 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1636968456
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1
transform 1 0 23828 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_263
timestamp 1636968456
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_275
timestamp 1
transform 1 0 25852 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_281
timestamp 1
transform 1 0 26404 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1
transform 1 0 28704 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_315
timestamp 1636968456
transform 1 0 29532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_327
timestamp 1
transform 1 0 30636 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636968456
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_27
timestamp 1
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_37
timestamp 1
transform 1 0 3956 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1
transform 1 0 4968 0 -1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636968456
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_69
timestamp 1
transform 1 0 6900 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_78
timestamp 1
transform 1 0 7728 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_86
timestamp 1
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_90
timestamp 1636968456
transform 1 0 8832 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_102
timestamp 1
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 1
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_140
timestamp 1636968456
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_152
timestamp 1
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_177
timestamp 1
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_191
timestamp 1
transform 1 0 18124 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_202
timestamp 1
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1
transform 1 0 20976 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_243
timestamp 1
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_263
timestamp 1636968456
transform 1 0 24748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_275
timestamp 1
transform 1 0 25852 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_291
timestamp 1636968456
transform 1 0 27324 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_303
timestamp 1
transform 1 0 28428 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_318
timestamp 1636968456
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_330
timestamp 1
transform 1 0 30912 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_334
timestamp 1
transform 1 0 31280 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636968456
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_55
timestamp 1636968456
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_67
timestamp 1
transform 1 0 6716 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_75
timestamp 1
transform 1 0 7452 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_115
timestamp 1
transform 1 0 11132 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_122
timestamp 1
transform 1 0 11776 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_130
timestamp 1
transform 1 0 12512 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1
transform 1 0 13524 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_166
timestamp 1
transform 1 0 15824 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_186
timestamp 1
transform 1 0 17664 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_215
timestamp 1636968456
transform 1 0 20332 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_227
timestamp 1
transform 1 0 21436 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_233
timestamp 1
transform 1 0 21988 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1
transform 1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636968456
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1636968456
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_277
timestamp 1
transform 1 0 26036 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_292
timestamp 1636968456
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_304
timestamp 1
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_318
timestamp 1636968456
transform 1 0 29808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_330
timestamp 1
transform 1 0 30912 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_334
timestamp 1
transform 1 0 31280 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 1
transform 1 0 1932 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_23
timestamp 1
transform 1 0 2668 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_38
timestamp 1
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_44
timestamp 1
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_63
timestamp 1
transform 1 0 6348 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_71
timestamp 1
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_89
timestamp 1
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_97
timestamp 1
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 1
transform 1 0 10028 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636968456
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636968456
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1636968456
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1636968456
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_180
timestamp 1
transform 1 0 17112 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_198
timestamp 1
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_206
timestamp 1
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_231
timestamp 1
transform 1 0 21804 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_239
timestamp 1
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_244
timestamp 1
transform 1 0 23000 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_248
timestamp 1
transform 1 0 23368 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_252
timestamp 1
transform 1 0 23736 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_261
timestamp 1
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_265
timestamp 1
transform 1 0 24932 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_269
timestamp 1
transform 1 0 25300 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1
transform 1 0 26036 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1636968456
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_305
timestamp 1
transform 1 0 28612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_318
timestamp 1636968456
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_330
timestamp 1
transform 1 0 30912 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_334
timestamp 1
transform 1 0 31280 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_15
timestamp 1
transform 1 0 1932 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_23
timestamp 1
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1
transform 1 0 3220 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_42
timestamp 1
transform 1 0 4416 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_57
timestamp 1
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_62
timestamp 1636968456
transform 1 0 6256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_74
timestamp 1
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_88
timestamp 1
transform 1 0 8648 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_129
timestamp 1
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_133
timestamp 1
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_146
timestamp 1
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_150
timestamp 1
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_154
timestamp 1636968456
transform 1 0 14720 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_166
timestamp 1
transform 1 0 15824 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 1
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_183
timestamp 1
transform 1 0 17388 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1636968456
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_209
timestamp 1
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_214
timestamp 1
transform 1 0 20240 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_220
timestamp 1
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_280
timestamp 1
transform 1 0 26312 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_295
timestamp 1
transform 1 0 27692 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_303
timestamp 1
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_318
timestamp 1636968456
transform 1 0 29808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_330
timestamp 1
transform 1 0 30912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_334
timestamp 1
transform 1 0 31280 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636968456
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_27
timestamp 1
transform 1 0 3036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1
transform 1 0 4140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_47
timestamp 1
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_87
timestamp 1
transform 1 0 8556 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_95
timestamp 1
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_107
timestamp 1
transform 1 0 10396 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636968456
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_146
timestamp 1
transform 1 0 13984 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_150
timestamp 1
transform 1 0 14352 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_163
timestamp 1
transform 1 0 15548 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_172
timestamp 1636968456
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_184
timestamp 1
transform 1 0 17480 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1636968456
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_237
timestamp 1
transform 1 0 22356 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_246
timestamp 1636968456
transform 1 0 23184 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_258
timestamp 1
transform 1 0 24288 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_266
timestamp 1
transform 1 0 25024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 1
transform 1 0 26404 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_289
timestamp 1
transform 1 0 27140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_303
timestamp 1
transform 1 0 28428 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1
transform 1 0 30820 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636968456
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636968456
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636968456
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp 1
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_64
timestamp 1636968456
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1
transform 1 0 8372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_93
timestamp 1
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_110
timestamp 1
transform 1 0 10672 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_114
timestamp 1
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_130
timestamp 1
transform 1 0 12512 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_150
timestamp 1
transform 1 0 14352 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_173
timestamp 1636968456
transform 1 0 16468 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_185
timestamp 1
transform 1 0 17572 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1636968456
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_209
timestamp 1
transform 1 0 19780 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_225
timestamp 1
transform 1 0 21252 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_233
timestamp 1
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1
transform 1 0 23552 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_268
timestamp 1
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_290
timestamp 1
transform 1 0 27232 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1
transform 1 0 28980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_317
timestamp 1
transform 1 0 29716 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_15
timestamp 1
transform 1 0 1932 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_23
timestamp 1
transform 1 0 2668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_36
timestamp 1
transform 1 0 3864 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_44
timestamp 1
transform 1 0 4600 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_92
timestamp 1
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_103
timestamp 1
transform 1 0 10028 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_126
timestamp 1636968456
transform 1 0 12144 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_147
timestamp 1
transform 1 0 14076 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_209
timestamp 1
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 1
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_225
timestamp 1
transform 1 0 21252 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_243
timestamp 1636968456
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_255
timestamp 1
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_269
timestamp 1
transform 1 0 25300 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1
transform 1 0 26036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_290
timestamp 1
transform 1 0 27232 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_298
timestamp 1
transform 1 0 27968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_309
timestamp 1
transform 1 0 28980 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_317
timestamp 1
transform 1 0 29716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_331
timestamp 1
transform 1 0 31004 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_15
timestamp 1
transform 1 0 1932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_32
timestamp 1
transform 1 0 3496 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_47
timestamp 1
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_54
timestamp 1
transform 1 0 5520 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_58
timestamp 1
transform 1 0 5888 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_62
timestamp 1636968456
transform 1 0 6256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636968456
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1636968456
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_109
timestamp 1
transform 1 0 10580 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_117
timestamp 1
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_127
timestamp 1
transform 1 0 12236 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_135
timestamp 1
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_147
timestamp 1
transform 1 0 14076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_155
timestamp 1
transform 1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_167
timestamp 1636968456
transform 1 0 15916 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_179
timestamp 1636968456
transform 1 0 17020 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 1
transform 1 0 18124 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_197
timestamp 1
transform 1 0 18676 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_218
timestamp 1
transform 1 0 20608 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_226
timestamp 1
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_240
timestamp 1636968456
transform 1 0 22632 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_253
timestamp 1
transform 1 0 23828 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_272
timestamp 1
transform 1 0 25576 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_276
timestamp 1
transform 1 0 25944 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_280
timestamp 1
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_291
timestamp 1
transform 1 0 27324 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_299
timestamp 1
transform 1 0 28060 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_306
timestamp 1
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_312
timestamp 1
transform 1 0 29256 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_330
timestamp 1
transform 1 0 30912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_334
timestamp 1
transform 1 0 31280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1
transform 1 0 828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_11
timestamp 1
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_28
timestamp 1
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_36
timestamp 1
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_49
timestamp 1
transform 1 0 5060 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_116
timestamp 1
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_133
timestamp 1
transform 1 0 12788 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_140
timestamp 1636968456
transform 1 0 13432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_152
timestamp 1
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_172
timestamp 1
transform 1 0 16376 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_180
timestamp 1
transform 1 0 17112 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_208
timestamp 1
transform 1 0 19688 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 1
transform 1 0 21252 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_243
timestamp 1636968456
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_255
timestamp 1
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_263
timestamp 1
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_270
timestamp 1
transform 1 0 25392 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1
transform 1 0 26036 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_284
timestamp 1636968456
transform 1 0 26680 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_296
timestamp 1
transform 1 0 27784 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_300
timestamp 1
transform 1 0 28152 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_313
timestamp 1
transform 1 0 29348 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_319
timestamp 1
transform 1 0 29900 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_24
timestamp 1
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_49
timestamp 1
transform 1 0 5060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp 1
transform 1 0 5612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_65
timestamp 1
transform 1 0 6532 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_72
timestamp 1636968456
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636968456
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_97
timestamp 1
transform 1 0 9476 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_105
timestamp 1
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_113
timestamp 1
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_119
timestamp 1
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_125
timestamp 1636968456
transform 1 0 12052 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636968456
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_153
timestamp 1
transform 1 0 14628 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_173
timestamp 1
transform 1 0 16468 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_179
timestamp 1
transform 1 0 17020 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_225
timestamp 1
transform 1 0 21252 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1
transform 1 0 23368 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1636968456
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_312
timestamp 1636968456
transform 1 0 29256 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_324
timestamp 1
transform 1 0 30360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_334
timestamp 1
transform 1 0 31280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_11
timestamp 1
transform 1 0 1564 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_27
timestamp 1
transform 1 0 3036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_35
timestamp 1
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_43
timestamp 1636968456
transform 1 0 4508 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_57
timestamp 1
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_66
timestamp 1
transform 1 0 6624 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_74
timestamp 1
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_100
timestamp 1
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_157
timestamp 1
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 1
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_176
timestamp 1
transform 1 0 16744 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_182
timestamp 1
transform 1 0 17296 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_198
timestamp 1636968456
transform 1 0 18768 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_210
timestamp 1
transform 1 0 19872 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1
transform 1 0 21252 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_245
timestamp 1
transform 1 0 23092 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_253
timestamp 1
transform 1 0 23828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_269
timestamp 1
transform 1 0 25300 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1
transform 1 0 26036 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636968456
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1636968456
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_305
timestamp 1
transform 1 0 28612 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_333
timestamp 1
transform 1 0 31188 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636968456
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_15
timestamp 1
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_32
timestamp 1
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_64
timestamp 1
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_69
timestamp 1
transform 1 0 6900 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_73
timestamp 1
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1
transform 1 0 8372 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1
transform 1 0 8924 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_98
timestamp 1636968456
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_113
timestamp 1
transform 1 0 10948 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_124
timestamp 1636968456
transform 1 0 11960 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp 1
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_158
timestamp 1636968456
transform 1 0 15088 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_170
timestamp 1
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_184
timestamp 1
transform 1 0 17480 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_192
timestamp 1
transform 1 0 18216 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_209
timestamp 1
transform 1 0 19780 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_213
timestamp 1
transform 1 0 20148 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_244
timestamp 1
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_264
timestamp 1636968456
transform 1 0 24840 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1636968456
transform 1 0 25944 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_288
timestamp 1636968456
transform 1 0 27048 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1
transform 1 0 28152 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_321
timestamp 1
transform 1 0 30084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_327
timestamp 1
transform 1 0 30636 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636968456
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_27
timestamp 1
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_35
timestamp 1
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_49
timestamp 1
transform 1 0 5060 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_61
timestamp 1
transform 1 0 6164 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_71
timestamp 1636968456
transform 1 0 7084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_83
timestamp 1
transform 1 0 8188 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_95
timestamp 1
transform 1 0 9292 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_99
timestamp 1
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_132
timestamp 1
transform 1 0 12696 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_142
timestamp 1
transform 1 0 13616 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_150
timestamp 1
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_169
timestamp 1
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_175
timestamp 1
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_188
timestamp 1
transform 1 0 17848 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_196
timestamp 1
transform 1 0 18584 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_211
timestamp 1636968456
transform 1 0 19964 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1
transform 1 0 21252 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_233
timestamp 1
transform 1 0 21988 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_237
timestamp 1
transform 1 0 22356 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1636968456
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1636968456
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1636968456
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_305
timestamp 1
transform 1 0 28612 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_323
timestamp 1636968456
transform 1 0 30268 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636968456
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_29
timestamp 1
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_50
timestamp 1
transform 1 0 5152 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_58
timestamp 1
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_101
timestamp 1636968456
transform 1 0 9844 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_113
timestamp 1
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_117
timestamp 1
transform 1 0 11316 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_124
timestamp 1
transform 1 0 11960 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_147
timestamp 1
transform 1 0 14076 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_153
timestamp 1
transform 1 0 14628 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_169
timestamp 1
transform 1 0 16100 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_175
timestamp 1
transform 1 0 16652 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_188
timestamp 1
transform 1 0 17848 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1
transform 1 0 18676 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_210
timestamp 1636968456
transform 1 0 19872 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_222
timestamp 1
transform 1 0 20976 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_230
timestamp 1
transform 1 0 21712 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_253
timestamp 1
transform 1 0 23828 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_259
timestamp 1
transform 1 0 24380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_271
timestamp 1
transform 1 0 25484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_327
timestamp 1
transform 1 0 30636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1
transform 1 0 828 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_11
timestamp 1
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_16
timestamp 1636968456
transform 1 0 2024 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_28
timestamp 1636968456
transform 1 0 3128 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_49
timestamp 1
transform 1 0 5060 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_66
timestamp 1
transform 1 0 6624 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_74
timestamp 1
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_85
timestamp 1
transform 1 0 8372 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_99
timestamp 1
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1
transform 1 0 10304 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_118
timestamp 1636968456
transform 1 0 11408 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_130
timestamp 1
transform 1 0 12512 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_136
timestamp 1
transform 1 0 13064 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_140
timestamp 1
transform 1 0 13432 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_150
timestamp 1
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_164
timestamp 1
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_169
timestamp 1
transform 1 0 16100 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_184
timestamp 1636968456
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_196
timestamp 1
transform 1 0 18584 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_209
timestamp 1
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_217
timestamp 1
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1
transform 1 0 20976 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_243
timestamp 1
transform 1 0 22908 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_251
timestamp 1
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_268
timestamp 1
transform 1 0 25208 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1636968456
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_293
timestamp 1
transform 1 0 27508 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_300
timestamp 1
transform 1 0 28152 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_308
timestamp 1
transform 1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_314
timestamp 1
transform 1 0 29440 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_320
timestamp 1636968456
transform 1 0 29992 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_332
timestamp 1
transform 1 0 31096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 1
transform 1 0 828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_32
timestamp 1
transform 1 0 3496 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_51
timestamp 1636968456
transform 1 0 5244 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_63
timestamp 1636968456
transform 1 0 6348 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_85
timestamp 1
transform 1 0 8372 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 1
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_150
timestamp 1
transform 1 0 14352 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_163
timestamp 1
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_177
timestamp 1
transform 1 0 16836 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_183
timestamp 1
transform 1 0 17388 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_206
timestamp 1
transform 1 0 19504 0 1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_226
timestamp 1636968456
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_238
timestamp 1
transform 1 0 22448 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_253
timestamp 1
transform 1 0 23828 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_266
timestamp 1636968456
transform 1 0 25024 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_278
timestamp 1
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_324
timestamp 1
transform 1 0 30360 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_332
timestamp 1
transform 1 0 31096 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 1
transform 1 0 828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_11
timestamp 1
transform 1 0 1564 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_24
timestamp 1
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_32
timestamp 1
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_47
timestamp 1
transform 1 0 4876 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_66
timestamp 1
transform 1 0 6624 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_79
timestamp 1
transform 1 0 7820 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_101
timestamp 1
transform 1 0 9844 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_109
timestamp 1
transform 1 0 10580 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636968456
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_125
timestamp 1
transform 1 0 12052 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_144
timestamp 1
transform 1 0 13800 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_152
timestamp 1
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636968456
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_181
timestamp 1
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_192
timestamp 1
transform 1 0 18216 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_203
timestamp 1
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1
transform 1 0 20792 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_225
timestamp 1
transform 1 0 21252 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_231
timestamp 1
transform 1 0 21804 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_271
timestamp 1
transform 1 0 25484 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_287
timestamp 1636968456
transform 1 0 26956 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_302
timestamp 1
transform 1 0 28336 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_310
timestamp 1
transform 1 0 29072 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_322
timestamp 1636968456
transform 1 0 30176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_334
timestamp 1
transform 1 0 31280 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_3
timestamp 1
transform 1 0 828 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_9
timestamp 1
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 1
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_43
timestamp 1636968456
transform 1 0 4508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_55
timestamp 1
transform 1 0 5612 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_68
timestamp 1
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_74
timestamp 1
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_85
timestamp 1
transform 1 0 8372 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_93
timestamp 1
transform 1 0 9108 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_112
timestamp 1636968456
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_124
timestamp 1
transform 1 0 11960 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_144
timestamp 1
transform 1 0 13800 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_164
timestamp 1
transform 1 0 15640 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_172
timestamp 1
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_202
timestamp 1
transform 1 0 19136 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_215
timestamp 1
transform 1 0 20332 0 1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_238
timestamp 1636968456
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1
transform 1 0 23552 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_253
timestamp 1
transform 1 0 23828 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_257
timestamp 1
transform 1 0 24196 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_264
timestamp 1
transform 1 0 24840 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_273
timestamp 1
transform 1 0 25668 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_280
timestamp 1636968456
transform 1 0 26312 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_292
timestamp 1
transform 1 0 27416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_300
timestamp 1
transform 1 0 28152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_304
timestamp 1
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1636968456
transform 1 0 30084 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_333
timestamp 1
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1
transform 1 0 828 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 1
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_22
timestamp 1
transform 1 0 2576 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_30
timestamp 1
transform 1 0 3312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_63
timestamp 1
transform 1 0 6348 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_86
timestamp 1
transform 1 0 8464 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_92
timestamp 1
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_99
timestamp 1
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_106
timestamp 1
transform 1 0 10304 0 -1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1636968456
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_140
timestamp 1
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_148
timestamp 1
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_189
timestamp 1
transform 1 0 17940 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_208
timestamp 1
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_234
timestamp 1636968456
transform 1 0 22080 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_276
timestamp 1
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1636968456
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_293
timestamp 1
transform 1 0 27508 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1636968456
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_321
timestamp 1636968456
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_333
timestamp 1
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_3
timestamp 1
transform 1 0 828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_9
timestamp 1
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_19
timestamp 1
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_23
timestamp 1
transform 1 0 2668 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_29
timestamp 1
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_33
timestamp 1
transform 1 0 3588 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_37
timestamp 1
transform 1 0 3956 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_44
timestamp 1
transform 1 0 4600 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_52
timestamp 1
transform 1 0 5336 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_56
timestamp 1636968456
transform 1 0 5704 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_68
timestamp 1
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_74
timestamp 1
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_88
timestamp 1
transform 1 0 8648 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_98
timestamp 1
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_106
timestamp 1
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_111
timestamp 1636968456
transform 1 0 10764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_123
timestamp 1
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_131
timestamp 1
transform 1 0 12604 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_144
timestamp 1
transform 1 0 13800 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_152
timestamp 1
transform 1 0 14536 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_158
timestamp 1
transform 1 0 15088 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_168
timestamp 1
transform 1 0 16008 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_176
timestamp 1
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_190
timestamp 1
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_206
timestamp 1
transform 1 0 19504 0 1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_224
timestamp 1636968456
transform 1 0 21160 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_236
timestamp 1
transform 1 0 22264 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1636968456
transform 1 0 23828 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_265
timestamp 1
transform 1 0 24932 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_274
timestamp 1
transform 1 0 25760 0 1 19040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1636968456
transform 1 0 26772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_297
timestamp 1
transform 1 0 27876 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_312
timestamp 1636968456
transform 1 0 29256 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_324
timestamp 1
transform 1 0 30360 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_332
timestamp 1
transform 1 0 31096 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_3
timestamp 1
transform 1 0 828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_62
timestamp 1
transform 1 0 6256 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_69
timestamp 1
transform 1 0 6900 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_77
timestamp 1
transform 1 0 7636 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_92
timestamp 1
transform 1 0 9016 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_101
timestamp 1
transform 1 0 9844 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_105
timestamp 1
transform 1 0 10212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_113
timestamp 1
transform 1 0 10948 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_126
timestamp 1
transform 1 0 12144 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_133
timestamp 1
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_153
timestamp 1
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_157
timestamp 1
transform 1 0 14996 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1
transform 1 0 15916 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_172
timestamp 1
transform 1 0 16376 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_178
timestamp 1
transform 1 0 16928 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_188
timestamp 1
transform 1 0 17848 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_194
timestamp 1
transform 1 0 18400 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_204
timestamp 1
transform 1 0 19320 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_219
timestamp 1
transform 1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_225
timestamp 1
transform 1 0 21252 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_248
timestamp 1
transform 1 0 23368 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_293
timestamp 1
transform 1 0 27508 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_299
timestamp 1
transform 1 0 28060 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_318
timestamp 1636968456
transform 1 0 29808 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_330
timestamp 1
transform 1 0 30912 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_334
timestamp 1
transform 1 0 31280 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1
transform 1 0 828 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_17
timestamp 1
transform 1 0 2116 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_25
timestamp 1
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_29
timestamp 1
transform 1 0 3220 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_38
timestamp 1636968456
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_50
timestamp 1636968456
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_62
timestamp 1
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_79
timestamp 1
transform 1 0 7820 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_88
timestamp 1636968456
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_100
timestamp 1636968456
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_112
timestamp 1
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_123
timestamp 1
transform 1 0 11868 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 1
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_149
timestamp 1
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_160
timestamp 1
transform 1 0 15272 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_174
timestamp 1
transform 1 0 16560 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_186
timestamp 1
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_192
timestamp 1
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_200
timestamp 1
transform 1 0 18952 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_212
timestamp 1
transform 1 0 20056 0 1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_229
timestamp 1636968456
transform 1 0 21620 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_241
timestamp 1
transform 1 0 22724 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_245
timestamp 1
transform 1 0 23092 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_262
timestamp 1636968456
transform 1 0 24656 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_274
timestamp 1
transform 1 0 25760 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_282
timestamp 1
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_295
timestamp 1636968456
transform 1 0 27692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_318
timestamp 1636968456
transform 1 0 29808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_330
timestamp 1
transform 1 0 30912 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_334
timestamp 1
transform 1 0 31280 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1636968456
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1636968456
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1636968456
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636968456
transform 1 0 5796 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1636968456
transform 1 0 6900 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1636968456
transform 1 0 8004 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1636968456
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1
transform 1 0 10212 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1636968456
transform 1 0 10948 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_125
timestamp 1
transform 1 0 12052 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_140
timestamp 1
transform 1 0 13432 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_144
timestamp 1
transform 1 0 13800 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_148
timestamp 1
transform 1 0 14168 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_152
timestamp 1
transform 1 0 14536 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 1
transform 1 0 15548 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_169
timestamp 1
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_187
timestamp 1
transform 1 0 17756 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_193
timestamp 1
transform 1 0 18308 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 1
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_252
timestamp 1
transform 1 0 23736 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_256
timestamp 1
transform 1 0 24104 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_264
timestamp 1
transform 1 0 24840 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_268
timestamp 1
transform 1 0 25208 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_276
timestamp 1
transform 1 0 25944 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_281
timestamp 1
transform 1 0 26404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_300
timestamp 1
transform 1 0 28152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_308
timestamp 1
transform 1 0 28888 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_321
timestamp 1636968456
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_333
timestamp 1
transform 1 0 31188 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1636968456
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636968456
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636968456
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_53
timestamp 1
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_57
timestamp 1
transform 1 0 5796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_64
timestamp 1
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_70
timestamp 1
transform 1 0 6992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_76
timestamp 1
transform 1 0 7544 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_88
timestamp 1
transform 1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_94
timestamp 1
transform 1 0 9200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_100
timestamp 1
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_106
timestamp 1
transform 1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_113
timestamp 1
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_118
timestamp 1
transform 1 0 11408 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_124
timestamp 1
transform 1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 1
transform 1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_136
timestamp 1
transform 1 0 13064 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_144
timestamp 1
transform 1 0 13800 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_148
timestamp 1
transform 1 0 14168 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_154
timestamp 1
transform 1 0 14720 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_167
timestamp 1
transform 1 0 15916 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_172
timestamp 1
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_181
timestamp 1
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_187
timestamp 1
transform 1 0 17756 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_191
timestamp 1
transform 1 0 18124 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_197
timestamp 1
transform 1 0 18676 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_203
timestamp 1
transform 1 0 19228 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_211
timestamp 1
transform 1 0 19964 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_244
timestamp 1
transform 1 0 23000 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_268
timestamp 1
transform 1 0 25208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_318
timestamp 1636968456
transform 1 0 29808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_330
timestamp 1
transform 1 0 30912 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_334
timestamp 1
transform 1 0 31280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 29532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 28612 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform 1 0 28428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform 1 0 27324 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform 1 0 27048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform 1 0 26036 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 26036 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 25208 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 24932 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform -1 0 23736 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform -1 0 23000 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform 1 0 22448 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform 1 0 22172 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform -1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1
transform -1 0 21528 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1
transform -1 0 20608 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1
transform -1 0 19964 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[0\].sky_inverter
timestamp 1
transform 1 0 20056 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[1\].sky_inverter
timestamp 1
transform 1 0 20332 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[2\].sky_inverter
timestamp 1
transform 1 0 20608 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[3\].sky_inverter
timestamp 1
transform 1 0 20792 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[4\].sky_inverter
timestamp 1
transform 1 0 21068 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[5\].sky_inverter
timestamp 1
transform 1 0 21344 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[6\].sky_inverter
timestamp 1
transform 1 0 21436 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[7\].sky_inverter
timestamp 1
transform 1 0 21712 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[8\].sky_inverter
timestamp 1
transform 1 0 21988 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[9\].sky_inverter
timestamp 1
transform 1 0 22264 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[10\].sky_inverter
timestamp 1
transform 1 0 22540 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[11\].sky_inverter
timestamp 1
transform 1 0 22816 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[12\].sky_inverter
timestamp 1
transform 1 0 23092 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[13\].sky_inverter
timestamp 1
transform -1 0 22908 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[14\].sky_inverter
timestamp 1
transform 1 0 23184 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[15\].sky_inverter
timestamp 1
transform -1 0 23184 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[16\].sky_inverter
timestamp 1
transform 1 0 23460 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[17\].sky_inverter
timestamp 1
transform -1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[18\].sky_inverter
timestamp 1
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[19\].sky_inverter
timestamp 1
transform 1 0 23736 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[20\].sky_inverter
timestamp 1
transform 1 0 24012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[21\].sky_inverter
timestamp 1
transform 1 0 24288 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[22\].sky_inverter
timestamp 1
transform 1 0 24564 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[23\].sky_inverter
timestamp 1
transform 1 0 24840 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[24\].sky_inverter
timestamp 1
transform 1 0 25116 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[25\].sky_inverter
timestamp 1
transform 1 0 25392 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[26\].sky_inverter
timestamp 1
transform 1 0 25668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[27\].sky_inverter
timestamp 1
transform -1 0 25668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[28\].sky_inverter
timestamp 1
transform 1 0 26036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[29\].sky_inverter
timestamp 1
transform -1 0 26036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[30\].sky_inverter
timestamp 1
transform 1 0 25760 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[31\].sky_inverter
timestamp 1
transform 1 0 26404 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[32\].sky_inverter
timestamp 1
transform 1 0 26680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[33\].sky_inverter
timestamp 1
transform -1 0 26312 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[34\].sky_inverter
timestamp 1
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[35\].sky_inverter
timestamp 1
transform 1 0 26588 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[36\].sky_inverter
timestamp 1
transform 1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[37\].sky_inverter
timestamp 1
transform 1 0 27140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[38\].sky_inverter
timestamp 1
transform 1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[39\].sky_inverter
timestamp 1
transform 1 0 27692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[40\].sky_inverter
timestamp 1
transform 1 0 27968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[41\].sky_inverter
timestamp 1
transform 1 0 28244 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[42\].sky_inverter
timestamp 1
transform 1 0 28520 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[43\].sky_inverter
timestamp 1
transform -1 0 28152 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[44\].sky_inverter
timestamp 1
transform 1 0 28060 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[45\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[46\].sky_inverter
timestamp 1
transform 1 0 29256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[47\].sky_inverter
timestamp 1
transform 1 0 29532 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[48\].sky_inverter
timestamp 1
transform 1 0 29808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[49\].sky_inverter
timestamp 1
transform -1 0 29440 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[50\].sky_inverter
timestamp 1
transform 1 0 30084 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[51\].sky_inverter
timestamp 1
transform -1 0 29624 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[52\].sky_inverter
timestamp 1
transform 1 0 29624 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[53\].sky_inverter
timestamp 1
transform 1 0 29900 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[54\].sky_inverter
timestamp 1
transform -1 0 29808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[55\].sky_inverter
timestamp 1
transform 1 0 29808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[56\].sky_inverter
timestamp 1
transform -1 0 29532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[57\].sky_inverter
timestamp 1
transform -1 0 29256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[58\].sky_inverter
timestamp 1
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[59\].sky_inverter
timestamp 1
transform 1 0 28704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[60\].sky_inverter
timestamp 1
transform -1 0 28520 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[61\].sky_inverter
timestamp 1
transform 1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[62\].sky_inverter
timestamp 1
transform -1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[63\].sky_inverter
timestamp 1
transform -1 0 28152 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[64\].sky_inverter
timestamp 1
transform 1 0 28060 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[65\].sky_inverter
timestamp 1
transform 1 0 28336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[66\].sky_inverter
timestamp 1
transform 1 0 28612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[67\].sky_inverter
timestamp 1
transform -1 0 28428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[68\].sky_inverter
timestamp 1
transform 1 0 28428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[69\].sky_inverter
timestamp 1
transform 1 0 28704 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[70\].sky_inverter
timestamp 1
transform 1 0 28980 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[71\].sky_inverter
timestamp 1
transform 1 0 29256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[72\].sky_inverter
timestamp 1
transform 1 0 29532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[73\].sky_inverter
timestamp 1
transform -1 0 29256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[74\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[75\].sky_inverter
timestamp 1
transform 1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[76\].sky_inverter
timestamp 1
transform 1 0 29532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[77\].sky_inverter
timestamp 1
transform -1 0 29256 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[78\].sky_inverter
timestamp 1
transform 1 0 29532 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[79\].sky_inverter
timestamp 1
transform 1 0 29808 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[80\].sky_inverter
timestamp 1
transform -1 0 29532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[81\].sky_inverter
timestamp 1
transform 1 0 29256 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[82\].sky_inverter
timestamp 1
transform -1 0 28612 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[83\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[84\].sky_inverter
timestamp 1
transform -1 0 28428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[85\].sky_inverter
timestamp 1
transform -1 0 28152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[86\].sky_inverter
timestamp 1
transform -1 0 27876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[87\].sky_inverter
timestamp 1
transform 1 0 27876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[88\].sky_inverter
timestamp 1
transform -1 0 27876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[89\].sky_inverter
timestamp 1
transform -1 0 27600 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[90\].sky_inverter
timestamp 1
transform -1 0 27324 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[91\].sky_inverter
timestamp 1
transform -1 0 27048 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[92\].sky_inverter
timestamp 1
transform 1 0 27416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[93\].sky_inverter
timestamp 1
transform -1 0 27416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[94\].sky_inverter
timestamp 1
transform -1 0 27140 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[95\].sky_inverter
timestamp 1
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[96\].sky_inverter
timestamp 1
transform -1 0 26772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[97\].sky_inverter
timestamp 1
transform 1 0 27232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[98\].sky_inverter
timestamp 1
transform -1 0 27232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[99\].sky_inverter
timestamp 1
transform -1 0 26956 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[100\].sky_inverter
timestamp 1
transform -1 0 26680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[101\].sky_inverter
timestamp 1
transform -1 0 25760 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[102\].sky_inverter
timestamp 1
transform 1 0 26036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[103\].sky_inverter
timestamp 1
transform -1 0 26036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[104\].sky_inverter
timestamp 1
transform -1 0 25760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[105\].sky_inverter
timestamp 1
transform -1 0 25484 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[106\].sky_inverter
timestamp 1
transform -1 0 25208 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[107\].sky_inverter
timestamp 1
transform -1 0 24932 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[108\].sky_inverter
timestamp 1
transform -1 0 24656 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[109\].sky_inverter
timestamp 1
transform -1 0 24380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[110\].sky_inverter
timestamp 1
transform 1 0 24380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[111\].sky_inverter
timestamp 1
transform -1 0 24380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[112\].sky_inverter
timestamp 1
transform -1 0 24104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[113\].sky_inverter
timestamp 1
transform -1 0 23736 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[114\].sky_inverter
timestamp 1
transform -1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[115\].sky_inverter
timestamp 1
transform -1 0 23460 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[116\].sky_inverter
timestamp 1
transform -1 0 23184 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[117\].sky_inverter
timestamp 1
transform -1 0 22908 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[118\].sky_inverter
timestamp 1
transform -1 0 22632 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[119\].sky_inverter
timestamp 1
transform -1 0 22356 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[120\].sky_inverter
timestamp 1
transform -1 0 22080 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[121\].sky_inverter
timestamp 1
transform -1 0 21528 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[122\].sky_inverter
timestamp 1
transform -1 0 21160 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[123\].sky_inverter
timestamp 1
transform -1 0 20884 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_62.inv_array\[124\].sky_inverter
timestamp 1
transform -1 0 20332 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[0\].sky_inverter
timestamp 1
transform -1 0 18952 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[1\].sky_inverter
timestamp 1
transform -1 0 18676 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[2\].sky_inverter
timestamp 1
transform -1 0 18584 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[3\].sky_inverter
timestamp 1
transform 1 0 18676 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[4\].sky_inverter
timestamp 1
transform 1 0 19044 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[5\].sky_inverter
timestamp 1
transform -1 0 19044 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[6\].sky_inverter
timestamp 1
transform -1 0 18768 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[7\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[8\].sky_inverter
timestamp 1
transform -1 0 19228 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[9\].sky_inverter
timestamp 1
transform -1 0 18952 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[10\].sky_inverter
timestamp 1
transform -1 0 18860 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[11\].sky_inverter
timestamp 1
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[12\].sky_inverter
timestamp 1
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[13\].sky_inverter
timestamp 1
transform -1 0 19136 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[14\].sky_inverter
timestamp 1
transform 1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[15\].sky_inverter
timestamp 1
transform 1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[16\].sky_inverter
timestamp 1
transform 1 0 19504 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[17\].sky_inverter
timestamp 1
transform 1 0 19780 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[18\].sky_inverter
timestamp 1
transform -1 0 19504 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[19\].sky_inverter
timestamp 1
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[20\].sky_inverter
timestamp 1
transform -1 0 19688 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[21\].sky_inverter
timestamp 1
transform 1 0 19688 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[22\].sky_inverter
timestamp 1
transform 1 0 19964 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[23\].sky_inverter
timestamp 1
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[24\].sky_inverter
timestamp 1
transform -1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[25\].sky_inverter
timestamp 1
transform 1 0 20240 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[26\].sky_inverter
timestamp 1
transform 1 0 20792 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[27\].sky_inverter
timestamp 1
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[28\].sky_inverter
timestamp 1
transform -1 0 20792 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[29\].sky_inverter
timestamp 1
transform 1 0 20700 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[30\].sky_inverter
timestamp 1
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[31\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[32\].sky_inverter
timestamp 1
transform 1 0 21804 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[33\].sky_inverter
timestamp 1
transform 1 0 22080 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[34\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[35\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[36\].sky_inverter
timestamp 1
transform -1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[37\].sky_inverter
timestamp 1
transform 1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[38\].sky_inverter
timestamp 1
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[39\].sky_inverter
timestamp 1
transform 1 0 22816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[40\].sky_inverter
timestamp 1
transform 1 0 23092 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[41\].sky_inverter
timestamp 1
transform 1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[42\].sky_inverter
timestamp 1
transform -1 0 23184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[43\].sky_inverter
timestamp 1
transform 1 0 23184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[44\].sky_inverter
timestamp 1
transform 1 0 23460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[45\].sky_inverter
timestamp 1
transform 1 0 24012 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[46\].sky_inverter
timestamp 1
transform -1 0 24012 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[47\].sky_inverter
timestamp 1
transform 1 0 24288 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[48\].sky_inverter
timestamp 1
transform -1 0 23736 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[49\].sky_inverter
timestamp 1
transform -1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[50\].sky_inverter
timestamp 1
transform 1 0 24288 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[51\].sky_inverter
timestamp 1
transform 1 0 24564 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[52\].sky_inverter
timestamp 1
transform -1 0 24288 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[53\].sky_inverter
timestamp 1
transform -1 0 24196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[54\].sky_inverter
timestamp 1
transform 1 0 24196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[55\].sky_inverter
timestamp 1
transform 1 0 24472 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[56\].sky_inverter
timestamp 1
transform 1 0 24748 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[57\].sky_inverter
timestamp 1
transform 1 0 25024 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[58\].sky_inverter
timestamp 1
transform -1 0 25208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[59\].sky_inverter
timestamp 1
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[60\].sky_inverter
timestamp 1
transform 1 0 25484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[61\].sky_inverter
timestamp 1
transform 1 0 25760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[62\].sky_inverter
timestamp 1
transform 1 0 26036 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[63\].sky_inverter
timestamp 1
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[64\].sky_inverter
timestamp 1
transform 1 0 26588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[65\].sky_inverter
timestamp 1
transform 1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[66\].sky_inverter
timestamp 1
transform 1 0 27140 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[67\].sky_inverter
timestamp 1
transform 1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[68\].sky_inverter
timestamp 1
transform 1 0 27692 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[69\].sky_inverter
timestamp 1
transform 1 0 27968 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[70\].sky_inverter
timestamp 1
transform 1 0 28244 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[71\].sky_inverter
timestamp 1
transform 1 0 28520 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[72\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[73\].sky_inverter
timestamp 1
transform 1 0 29072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[74\].sky_inverter
timestamp 1
transform -1 0 29072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[75\].sky_inverter
timestamp 1
transform -1 0 28796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[76\].sky_inverter
timestamp 1
transform -1 0 28520 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[77\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[78\].sky_inverter
timestamp 1
transform -1 0 28704 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[79\].sky_inverter
timestamp 1
transform -1 0 28428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[80\].sky_inverter
timestamp 1
transform 1 0 28704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[81\].sky_inverter
timestamp 1
transform -1 0 28704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[82\].sky_inverter
timestamp 1
transform -1 0 28428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[83\].sky_inverter
timestamp 1
transform -1 0 28336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[84\].sky_inverter
timestamp 1
transform 1 0 28336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[85\].sky_inverter
timestamp 1
transform 1 0 28612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[86\].sky_inverter
timestamp 1
transform -1 0 28060 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[87\].sky_inverter
timestamp 1
transform 1 0 28152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[88\].sky_inverter
timestamp 1
transform -1 0 28152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[89\].sky_inverter
timestamp 1
transform -1 0 27876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[90\].sky_inverter
timestamp 1
transform -1 0 27600 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[91\].sky_inverter
timestamp 1
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[92\].sky_inverter
timestamp 1
transform 1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[93\].sky_inverter
timestamp 1
transform -1 0 27140 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[94\].sky_inverter
timestamp 1
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[95\].sky_inverter
timestamp 1
transform 1 0 26680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[96\].sky_inverter
timestamp 1
transform 1 0 26956 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[97\].sky_inverter
timestamp 1
transform 1 0 27232 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[98\].sky_inverter
timestamp 1
transform -1 0 26680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[99\].sky_inverter
timestamp 1
transform 1 0 26588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[100\].sky_inverter
timestamp 1
transform 1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[101\].sky_inverter
timestamp 1
transform 1 0 27140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[102\].sky_inverter
timestamp 1
transform -1 0 26588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[103\].sky_inverter
timestamp 1
transform 1 0 26496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[104\].sky_inverter
timestamp 1
transform 1 0 26772 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[105\].sky_inverter
timestamp 1
transform 1 0 27048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[106\].sky_inverter
timestamp 1
transform -1 0 26772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[107\].sky_inverter
timestamp 1
transform 1 0 26772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[108\].sky_inverter
timestamp 1
transform 1 0 27048 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[109\].sky_inverter
timestamp 1
transform 1 0 27324 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[110\].sky_inverter
timestamp 1
transform 1 0 27600 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[111\].sky_inverter
timestamp 1
transform 1 0 27876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[112\].sky_inverter
timestamp 1
transform 1 0 28152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[113\].sky_inverter
timestamp 1
transform 1 0 28428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[114\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[115\].sky_inverter
timestamp 1
transform -1 0 29164 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[116\].sky_inverter
timestamp 1
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[117\].sky_inverter
timestamp 1
transform 1 0 29256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[118\].sky_inverter
timestamp 1
transform 1 0 29532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[119\].sky_inverter
timestamp 1
transform -1 0 29532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[120\].sky_inverter
timestamp 1
transform -1 0 29256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[121\].sky_inverter
timestamp 1
transform -1 0 28980 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[122\].sky_inverter
timestamp 1
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[123\].sky_inverter
timestamp 1
transform 1 0 29532 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[124\].sky_inverter
timestamp 1
transform -1 0 29532 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[125\].sky_inverter
timestamp 1
transform -1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[126\].sky_inverter
timestamp 1
transform 1 0 29532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[127\].sky_inverter
timestamp 1
transform -1 0 29532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[128\].sky_inverter
timestamp 1
transform -1 0 29256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[129\].sky_inverter
timestamp 1
transform -1 0 28980 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[130\].sky_inverter
timestamp 1
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[131\].sky_inverter
timestamp 1
transform 1 0 29532 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[132\].sky_inverter
timestamp 1
transform -1 0 29256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[133\].sky_inverter
timestamp 1
transform 1 0 29256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[134\].sky_inverter
timestamp 1
transform -1 0 29440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[135\].sky_inverter
timestamp 1
transform 1 0 29440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[136\].sky_inverter
timestamp 1
transform 1 0 29716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[137\].sky_inverter
timestamp 1
transform 1 0 29992 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[138\].sky_inverter
timestamp 1
transform 1 0 30268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[139\].sky_inverter
timestamp 1
transform 1 0 30544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[140\].sky_inverter
timestamp 1
transform -1 0 30268 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[141\].sky_inverter
timestamp 1
transform 1 0 31096 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[142\].sky_inverter
timestamp 1
transform -1 0 31096 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[143\].sky_inverter
timestamp 1
transform -1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[144\].sky_inverter
timestamp 1
transform -1 0 30544 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[145\].sky_inverter
timestamp 1
transform -1 0 30452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[146\].sky_inverter
timestamp 1
transform 1 0 30452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[147\].sky_inverter
timestamp 1
transform -1 0 30176 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[148\].sky_inverter
timestamp 1
transform 1 0 30728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[149\].sky_inverter
timestamp 1
transform -1 0 30084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[150\].sky_inverter
timestamp 1
transform 1 0 30084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[151\].sky_inverter
timestamp 1
transform 1 0 30360 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[152\].sky_inverter
timestamp 1
transform 1 0 30636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[153\].sky_inverter
timestamp 1
transform -1 0 30268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[154\].sky_inverter
timestamp 1
transform 1 0 30268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[155\].sky_inverter
timestamp 1
transform 1 0 30544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[156\].sky_inverter
timestamp 1
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[157\].sky_inverter
timestamp 1
transform 1 0 31096 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[158\].sky_inverter
timestamp 1
transform -1 0 30728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[159\].sky_inverter
timestamp 1
transform 1 0 30728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[160\].sky_inverter
timestamp 1
transform 1 0 31004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[161\].sky_inverter
timestamp 1
transform -1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[162\].sky_inverter
timestamp 1
transform 1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[163\].sky_inverter
timestamp 1
transform -1 0 30636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[164\].sky_inverter
timestamp 1
transform 1 0 30360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[165\].sky_inverter
timestamp 1
transform -1 0 30360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[166\].sky_inverter
timestamp 1
transform -1 0 30084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[167\].sky_inverter
timestamp 1
transform -1 0 29808 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[168\].sky_inverter
timestamp 1
transform -1 0 29532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[169\].sky_inverter
timestamp 1
transform -1 0 29256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[170\].sky_inverter
timestamp 1
transform 1 0 28980 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[171\].sky_inverter
timestamp 1
transform 1 0 29256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[172\].sky_inverter
timestamp 1
transform 1 0 29532 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[173\].sky_inverter
timestamp 1
transform 1 0 29808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[174\].sky_inverter
timestamp 1
transform -1 0 29440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[175\].sky_inverter
timestamp 1
transform 1 0 29440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[176\].sky_inverter
timestamp 1
transform 1 0 29716 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[177\].sky_inverter
timestamp 1
transform 1 0 29992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[178\].sky_inverter
timestamp 1
transform 1 0 30084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[179\].sky_inverter
timestamp 1
transform -1 0 29992 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[180\].sky_inverter
timestamp 1
transform 1 0 30360 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[181\].sky_inverter
timestamp 1
transform -1 0 30084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[182\].sky_inverter
timestamp 1
transform -1 0 29808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[183\].sky_inverter
timestamp 1
transform -1 0 29532 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[184\].sky_inverter
timestamp 1
transform -1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[185\].sky_inverter
timestamp 1
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[186\].sky_inverter
timestamp 1
transform -1 0 28612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[187\].sky_inverter
timestamp 1
transform -1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[188\].sky_inverter
timestamp 1
transform -1 0 28060 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[189\].sky_inverter
timestamp 1
transform -1 0 27784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[190\].sky_inverter
timestamp 1
transform -1 0 27508 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[191\].sky_inverter
timestamp 1
transform -1 0 27232 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[192\].sky_inverter
timestamp 1
transform -1 0 26956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[193\].sky_inverter
timestamp 1
transform -1 0 26680 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[194\].sky_inverter
timestamp 1
transform -1 0 26404 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[195\].sky_inverter
timestamp 1
transform -1 0 26128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[196\].sky_inverter
timestamp 1
transform -1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[197\].sky_inverter
timestamp 1
transform -1 0 25852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[198\].sky_inverter
timestamp 1
transform -1 0 25576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[199\].sky_inverter
timestamp 1
transform -1 0 25484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[200\].sky_inverter
timestamp 1
transform -1 0 25208 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[201\].sky_inverter
timestamp 1
transform -1 0 24932 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[202\].sky_inverter
timestamp 1
transform 1 0 24932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[203\].sky_inverter
timestamp 1
transform -1 0 24932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[204\].sky_inverter
timestamp 1
transform -1 0 24380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[205\].sky_inverter
timestamp 1
transform 1 0 24380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[206\].sky_inverter
timestamp 1
transform -1 0 24104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[207\].sky_inverter
timestamp 1
transform 1 0 24104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[208\].sky_inverter
timestamp 1
transform 1 0 24196 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[209\].sky_inverter
timestamp 1
transform 1 0 24472 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[210\].sky_inverter
timestamp 1
transform 1 0 24748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[211\].sky_inverter
timestamp 1
transform 1 0 25208 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[212\].sky_inverter
timestamp 1
transform -1 0 24840 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[213\].sky_inverter
timestamp 1
transform -1 0 24564 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[214\].sky_inverter
timestamp 1
transform 1 0 24932 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[215\].sky_inverter
timestamp 1
transform -1 0 24932 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[216\].sky_inverter
timestamp 1
transform -1 0 24656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[217\].sky_inverter
timestamp 1
transform -1 0 24380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[218\].sky_inverter
timestamp 1
transform -1 0 24104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[219\].sky_inverter
timestamp 1
transform -1 0 23092 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[220\].sky_inverter
timestamp 1
transform 1 0 23552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[221\].sky_inverter
timestamp 1
transform -1 0 23552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[222\].sky_inverter
timestamp 1
transform -1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[223\].sky_inverter
timestamp 1
transform -1 0 23000 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[224\].sky_inverter
timestamp 1
transform -1 0 22724 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[225\].sky_inverter
timestamp 1
transform -1 0 22172 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[226\].sky_inverter
timestamp 1
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[227\].sky_inverter
timestamp 1
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[228\].sky_inverter
timestamp 1
transform 1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[229\].sky_inverter
timestamp 1
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[230\].sky_inverter
timestamp 1
transform 1 0 22172 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[231\].sky_inverter
timestamp 1
transform -1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[232\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[233\].sky_inverter
timestamp 1
transform 1 0 21804 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[234\].sky_inverter
timestamp 1
transform -1 0 20700 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[235\].sky_inverter
timestamp 1
transform 1 0 21252 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[236\].sky_inverter
timestamp 1
transform -1 0 20976 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[237\].sky_inverter
timestamp 1
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[238\].sky_inverter
timestamp 1
transform 1 0 20884 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[239\].sky_inverter
timestamp 1
transform -1 0 20608 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[240\].sky_inverter
timestamp 1
transform -1 0 20332 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[241\].sky_inverter
timestamp 1
transform 1 0 20148 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[242\].sky_inverter
timestamp 1
transform 1 0 20424 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[243\].sky_inverter
timestamp 1
transform -1 0 20148 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[244\].sky_inverter
timestamp 1
transform -1 0 19872 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[245\].sky_inverter
timestamp 1
transform -1 0 19780 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[246\].sky_inverter
timestamp 1
transform 1 0 19780 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[247\].sky_inverter
timestamp 1
transform -1 0 20056 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[248\].sky_inverter
timestamp 1
transform -1 0 19780 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[249\].sky_inverter
timestamp 1
transform -1 0 19504 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_125.inv_array\[250\].sky_inverter
timestamp 1
transform -1 0 19228 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[0\].sky_inverter
timestamp 1
transform -1 0 17480 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[1\].sky_inverter
timestamp 1
transform -1 0 17204 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[2\].sky_inverter
timestamp 1
transform -1 0 16928 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[3\].sky_inverter
timestamp 1
transform -1 0 16652 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[4\].sky_inverter
timestamp 1
transform -1 0 16560 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[5\].sky_inverter
timestamp 1
transform -1 0 16284 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[6\].sky_inverter
timestamp 1
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[7\].sky_inverter
timestamp 1
transform -1 0 15916 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[8\].sky_inverter
timestamp 1
transform -1 0 15640 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[9\].sky_inverter
timestamp 1
transform -1 0 15364 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[10\].sky_inverter
timestamp 1
transform 1 0 15180 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[11\].sky_inverter
timestamp 1
transform 1 0 15732 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[12\].sky_inverter
timestamp 1
transform -1 0 15732 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[13\].sky_inverter
timestamp 1
transform -1 0 15088 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[14\].sky_inverter
timestamp 1
transform -1 0 14720 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[15\].sky_inverter
timestamp 1
transform 1 0 15548 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[16\].sky_inverter
timestamp 1
transform -1 0 15548 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[17\].sky_inverter
timestamp 1
transform -1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[18\].sky_inverter
timestamp 1
transform -1 0 14996 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[19\].sky_inverter
timestamp 1
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[20\].sky_inverter
timestamp 1
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[21\].sky_inverter
timestamp 1
transform -1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[22\].sky_inverter
timestamp 1
transform -1 0 15088 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[23\].sky_inverter
timestamp 1
transform -1 0 14996 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[24\].sky_inverter
timestamp 1
transform 1 0 15548 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[25\].sky_inverter
timestamp 1
transform -1 0 15548 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[26\].sky_inverter
timestamp 1
transform -1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[27\].sky_inverter
timestamp 1
transform 1 0 14996 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[28\].sky_inverter
timestamp 1
transform 1 0 15364 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[29\].sky_inverter
timestamp 1
transform -1 0 15364 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[30\].sky_inverter
timestamp 1
transform -1 0 14996 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[31\].sky_inverter
timestamp 1
transform 1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[32\].sky_inverter
timestamp 1
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[33\].sky_inverter
timestamp 1
transform -1 0 15548 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[34\].sky_inverter
timestamp 1
transform -1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[35\].sky_inverter
timestamp 1
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[36\].sky_inverter
timestamp 1
transform -1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[37\].sky_inverter
timestamp 1
transform -1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[38\].sky_inverter
timestamp 1
transform -1 0 15180 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[39\].sky_inverter
timestamp 1
transform -1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[40\].sky_inverter
timestamp 1
transform 1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[41\].sky_inverter
timestamp 1
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[42\].sky_inverter
timestamp 1
transform -1 0 14536 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[43\].sky_inverter
timestamp 1
transform -1 0 14444 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[44\].sky_inverter
timestamp 1
transform 1 0 14444 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[45\].sky_inverter
timestamp 1
transform 1 0 14720 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[46\].sky_inverter
timestamp 1
transform -1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[47\].sky_inverter
timestamp 1
transform -1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[48\].sky_inverter
timestamp 1
transform -1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[49\].sky_inverter
timestamp 1
transform -1 0 13340 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[50\].sky_inverter
timestamp 1
transform -1 0 13064 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[51\].sky_inverter
timestamp 1
transform -1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[52\].sky_inverter
timestamp 1
transform -1 0 12512 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[53\].sky_inverter
timestamp 1
transform -1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[54\].sky_inverter
timestamp 1
transform -1 0 11960 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[55\].sky_inverter
timestamp 1
transform -1 0 11684 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[56\].sky_inverter
timestamp 1
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[57\].sky_inverter
timestamp 1
transform -1 0 11408 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[58\].sky_inverter
timestamp 1
transform 1 0 11224 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[59\].sky_inverter
timestamp 1
transform -1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[60\].sky_inverter
timestamp 1
transform -1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[61\].sky_inverter
timestamp 1
transform 1 0 10672 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[62\].sky_inverter
timestamp 1
transform -1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[63\].sky_inverter
timestamp 1
transform -1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[64\].sky_inverter
timestamp 1
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[65\].sky_inverter
timestamp 1
transform -1 0 10672 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[66\].sky_inverter
timestamp 1
transform -1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[67\].sky_inverter
timestamp 1
transform -1 0 10120 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[68\].sky_inverter
timestamp 1
transform -1 0 9844 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[69\].sky_inverter
timestamp 1
transform -1 0 9568 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[70\].sky_inverter
timestamp 1
transform -1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[71\].sky_inverter
timestamp 1
transform -1 0 9016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[72\].sky_inverter
timestamp 1
transform -1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[73\].sky_inverter
timestamp 1
transform -1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[74\].sky_inverter
timestamp 1
transform -1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[75\].sky_inverter
timestamp 1
transform -1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[76\].sky_inverter
timestamp 1
transform -1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[77\].sky_inverter
timestamp 1
transform -1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[78\].sky_inverter
timestamp 1
transform 1 0 7360 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[79\].sky_inverter
timestamp 1
transform -1 0 7084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[80\].sky_inverter
timestamp 1
transform -1 0 6808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[81\].sky_inverter
timestamp 1
transform 1 0 6624 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[82\].sky_inverter
timestamp 1
transform 1 0 6900 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[83\].sky_inverter
timestamp 1
transform -1 0 6532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[84\].sky_inverter
timestamp 1
transform -1 0 6256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[85\].sky_inverter
timestamp 1
transform -1 0 5980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[86\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[87\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[88\].sky_inverter
timestamp 1
transform 1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[89\].sky_inverter
timestamp 1
transform -1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[90\].sky_inverter
timestamp 1
transform -1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[91\].sky_inverter
timestamp 1
transform 1 0 6256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[92\].sky_inverter
timestamp 1
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[93\].sky_inverter
timestamp 1
transform 1 0 6808 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[94\].sky_inverter
timestamp 1
transform -1 0 6624 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[95\].sky_inverter
timestamp 1
transform 1 0 6624 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[96\].sky_inverter
timestamp 1
transform 1 0 6900 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[97\].sky_inverter
timestamp 1
transform -1 0 6348 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[98\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[99\].sky_inverter
timestamp 1
transform 1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[100\].sky_inverter
timestamp 1
transform -1 0 6072 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[101\].sky_inverter
timestamp 1
transform -1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[102\].sky_inverter
timestamp 1
transform -1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[103\].sky_inverter
timestamp 1
transform -1 0 5244 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[104\].sky_inverter
timestamp 1
transform -1 0 4692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[105\].sky_inverter
timestamp 1
transform -1 0 3864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[106\].sky_inverter
timestamp 1
transform -1 0 3496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[107\].sky_inverter
timestamp 1
transform -1 0 3036 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[108\].sky_inverter
timestamp 1
transform -1 0 2760 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[109\].sky_inverter
timestamp 1
transform -1 0 2484 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[110\].sky_inverter
timestamp 1
transform -1 0 2208 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[111\].sky_inverter
timestamp 1
transform -1 0 1932 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[112\].sky_inverter
timestamp 1
transform -1 0 1656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[113\].sky_inverter
timestamp 1
transform 1 0 1748 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[114\].sky_inverter
timestamp 1
transform -1 0 1932 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[115\].sky_inverter
timestamp 1
transform -1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[116\].sky_inverter
timestamp 1
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[117\].sky_inverter
timestamp 1
transform 1 0 2208 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[118\].sky_inverter
timestamp 1
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[119\].sky_inverter
timestamp 1
transform -1 0 2024 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[120\].sky_inverter
timestamp 1
transform 1 0 2024 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[121\].sky_inverter
timestamp 1
transform 1 0 2300 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[122\].sky_inverter
timestamp 1
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[123\].sky_inverter
timestamp 1
transform -1 0 1748 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[124\].sky_inverter
timestamp 1
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[125\].sky_inverter
timestamp 1
transform 1 0 2024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[126\].sky_inverter
timestamp 1
transform 1 0 2300 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[127\].sky_inverter
timestamp 1
transform -1 0 1748 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[128\].sky_inverter
timestamp 1
transform 1 0 1472 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[129\].sky_inverter
timestamp 1
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[130\].sky_inverter
timestamp 1
transform 1 0 2024 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[131\].sky_inverter
timestamp 1
transform -1 0 1564 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[132\].sky_inverter
timestamp 1
transform 1 0 1564 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[133\].sky_inverter
timestamp 1
transform -1 0 1288 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[134\].sky_inverter
timestamp 1
transform 1 0 1840 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[135\].sky_inverter
timestamp 1
transform -1 0 1840 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[136\].sky_inverter
timestamp 1
transform 1 0 1840 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[137\].sky_inverter
timestamp 1
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[138\].sky_inverter
timestamp 1
transform 1 0 2760 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[139\].sky_inverter
timestamp 1
transform -1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[140\].sky_inverter
timestamp 1
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[141\].sky_inverter
timestamp 1
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[142\].sky_inverter
timestamp 1
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[143\].sky_inverter
timestamp 1
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[144\].sky_inverter
timestamp 1
transform -1 0 3772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[145\].sky_inverter
timestamp 1
transform 1 0 3772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[146\].sky_inverter
timestamp 1
transform 1 0 4324 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[147\].sky_inverter
timestamp 1
transform -1 0 4324 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[148\].sky_inverter
timestamp 1
transform 1 0 4324 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[149\].sky_inverter
timestamp 1
transform 1 0 4600 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[150\].sky_inverter
timestamp 1
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[151\].sky_inverter
timestamp 1
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[152\].sky_inverter
timestamp 1
transform -1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[153\].sky_inverter
timestamp 1
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[154\].sky_inverter
timestamp 1
transform 1 0 5980 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[155\].sky_inverter
timestamp 1
transform 1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[156\].sky_inverter
timestamp 1
transform -1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[157\].sky_inverter
timestamp 1
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[158\].sky_inverter
timestamp 1
transform 1 0 6716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[159\].sky_inverter
timestamp 1
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[160\].sky_inverter
timestamp 1
transform 1 0 7268 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[161\].sky_inverter
timestamp 1
transform 1 0 7544 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[162\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[163\].sky_inverter
timestamp 1
transform -1 0 8188 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[164\].sky_inverter
timestamp 1
transform 1 0 8740 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[165\].sky_inverter
timestamp 1
transform -1 0 8740 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[166\].sky_inverter
timestamp 1
transform -1 0 8464 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[167\].sky_inverter
timestamp 1
transform -1 0 8188 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[168\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[169\].sky_inverter
timestamp 1
transform -1 0 8280 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[170\].sky_inverter
timestamp 1
transform -1 0 8004 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[171\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[172\].sky_inverter
timestamp 1
transform -1 0 7360 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[173\].sky_inverter
timestamp 1
transform 1 0 8188 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[174\].sky_inverter
timestamp 1
transform -1 0 8188 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[175\].sky_inverter
timestamp 1
transform -1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[176\].sky_inverter
timestamp 1
transform -1 0 7636 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[177\].sky_inverter
timestamp 1
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[178\].sky_inverter
timestamp 1
transform -1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[179\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[180\].sky_inverter
timestamp 1
transform -1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[181\].sky_inverter
timestamp 1
transform 1 0 7728 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[182\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[183\].sky_inverter
timestamp 1
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[184\].sky_inverter
timestamp 1
transform -1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[185\].sky_inverter
timestamp 1
transform -1 0 7820 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[186\].sky_inverter
timestamp 1
transform -1 0 7452 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[187\].sky_inverter
timestamp 1
transform 1 0 7452 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[188\].sky_inverter
timestamp 1
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[189\].sky_inverter
timestamp 1
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[190\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[191\].sky_inverter
timestamp 1
transform 1 0 8648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[192\].sky_inverter
timestamp 1
transform 1 0 9292 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[193\].sky_inverter
timestamp 1
transform 1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[194\].sky_inverter
timestamp 1
transform 1 0 9752 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[195\].sky_inverter
timestamp 1
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[196\].sky_inverter
timestamp 1
transform 1 0 10304 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[197\].sky_inverter
timestamp 1
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[198\].sky_inverter
timestamp 1
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[199\].sky_inverter
timestamp 1
transform -1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[200\].sky_inverter
timestamp 1
transform 1 0 11040 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[201\].sky_inverter
timestamp 1
transform 1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[202\].sky_inverter
timestamp 1
transform -1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[203\].sky_inverter
timestamp 1
transform 1 0 11592 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[204\].sky_inverter
timestamp 1
transform 1 0 11868 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[205\].sky_inverter
timestamp 1
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[206\].sky_inverter
timestamp 1
transform 1 0 12420 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[207\].sky_inverter
timestamp 1
transform 1 0 13340 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[208\].sky_inverter
timestamp 1
transform -1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[209\].sky_inverter
timestamp 1
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[210\].sky_inverter
timestamp 1
transform -1 0 13248 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[211\].sky_inverter
timestamp 1
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[212\].sky_inverter
timestamp 1
transform 1 0 13800 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[213\].sky_inverter
timestamp 1
transform -1 0 12972 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[214\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[215\].sky_inverter
timestamp 1
transform 1 0 14076 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[216\].sky_inverter
timestamp 1
transform -1 0 14076 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[217\].sky_inverter
timestamp 1
transform -1 0 13800 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[218\].sky_inverter
timestamp 1
transform 1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[219\].sky_inverter
timestamp 1
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[220\].sky_inverter
timestamp 1
transform 1 0 14444 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[221\].sky_inverter
timestamp 1
transform 1 0 14720 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[222\].sky_inverter
timestamp 1
transform 1 0 15272 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[223\].sky_inverter
timestamp 1
transform 1 0 15732 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[224\].sky_inverter
timestamp 1
transform 1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[225\].sky_inverter
timestamp 1
transform 1 0 16284 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[226\].sky_inverter
timestamp 1
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[227\].sky_inverter
timestamp 1
transform 1 0 16652 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[228\].sky_inverter
timestamp 1
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[229\].sky_inverter
timestamp 1
transform -1 0 17204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[230\].sky_inverter
timestamp 1
transform -1 0 17020 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[231\].sky_inverter
timestamp 1
transform 1 0 17572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[232\].sky_inverter
timestamp 1
transform -1 0 17572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[233\].sky_inverter
timestamp 1
transform -1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[234\].sky_inverter
timestamp 1
transform 1 0 17572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[235\].sky_inverter
timestamp 1
transform -1 0 17572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[236\].sky_inverter
timestamp 1
transform -1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[237\].sky_inverter
timestamp 1
transform -1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[238\].sky_inverter
timestamp 1
transform 1 0 17204 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[239\].sky_inverter
timestamp 1
transform -1 0 17204 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[240\].sky_inverter
timestamp 1
transform -1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[241\].sky_inverter
timestamp 1
transform -1 0 16652 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[242\].sky_inverter
timestamp 1
transform -1 0 16468 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[243\].sky_inverter
timestamp 1
transform 1 0 16468 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[244\].sky_inverter
timestamp 1
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[245\].sky_inverter
timestamp 1
transform -1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[246\].sky_inverter
timestamp 1
transform -1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[247\].sky_inverter
timestamp 1
transform 1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[248\].sky_inverter
timestamp 1
transform -1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[249\].sky_inverter
timestamp 1
transform -1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[250\].sky_inverter
timestamp 1
transform -1 0 15640 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[251\].sky_inverter
timestamp 1
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[252\].sky_inverter
timestamp 1
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[253\].sky_inverter
timestamp 1
transform -1 0 15916 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[254\].sky_inverter
timestamp 1
transform -1 0 15640 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[255\].sky_inverter
timestamp 1
transform 1 0 15640 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[256\].sky_inverter
timestamp 1
transform -1 0 15640 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[257\].sky_inverter
timestamp 1
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[258\].sky_inverter
timestamp 1
transform -1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[259\].sky_inverter
timestamp 1
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[260\].sky_inverter
timestamp 1
transform -1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[261\].sky_inverter
timestamp 1
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[262\].sky_inverter
timestamp 1
transform 1 0 15088 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[263\].sky_inverter
timestamp 1
transform 1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[264\].sky_inverter
timestamp 1
transform 1 0 15640 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[265\].sky_inverter
timestamp 1
transform 1 0 15916 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[266\].sky_inverter
timestamp 1
transform 1 0 16192 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[267\].sky_inverter
timestamp 1
transform 1 0 16468 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[268\].sky_inverter
timestamp 1
transform 1 0 16744 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[269\].sky_inverter
timestamp 1
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[270\].sky_inverter
timestamp 1
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[271\].sky_inverter
timestamp 1
transform 1 0 17572 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[272\].sky_inverter
timestamp 1
transform 1 0 17848 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[273\].sky_inverter
timestamp 1
transform 1 0 18124 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[274\].sky_inverter
timestamp 1
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[275\].sky_inverter
timestamp 1
transform 1 0 18676 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[276\].sky_inverter
timestamp 1
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[277\].sky_inverter
timestamp 1
transform 1 0 19228 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[278\].sky_inverter
timestamp 1
transform 1 0 19504 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[279\].sky_inverter
timestamp 1
transform -1 0 19228 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[280\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[281\].sky_inverter
timestamp 1
transform 1 0 19504 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[282\].sky_inverter
timestamp 1
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[283\].sky_inverter
timestamp 1
transform 1 0 20056 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[284\].sky_inverter
timestamp 1
transform 1 0 20332 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[285\].sky_inverter
timestamp 1
transform -1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[286\].sky_inverter
timestamp 1
transform 1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[287\].sky_inverter
timestamp 1
transform -1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[288\].sky_inverter
timestamp 1
transform 1 0 20424 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[289\].sky_inverter
timestamp 1
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[290\].sky_inverter
timestamp 1
transform 1 0 20976 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[291\].sky_inverter
timestamp 1
transform -1 0 20424 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[292\].sky_inverter
timestamp 1
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[293\].sky_inverter
timestamp 1
transform -1 0 20240 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[294\].sky_inverter
timestamp 1
transform 1 0 20608 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[295\].sky_inverter
timestamp 1
transform -1 0 20608 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[296\].sky_inverter
timestamp 1
transform -1 0 20332 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[297\].sky_inverter
timestamp 1
transform -1 0 20056 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[298\].sky_inverter
timestamp 1
transform -1 0 19780 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[299\].sky_inverter
timestamp 1
transform -1 0 19504 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[300\].sky_inverter
timestamp 1
transform -1 0 19228 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[301\].sky_inverter
timestamp 1
transform -1 0 18952 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[302\].sky_inverter
timestamp 1
transform -1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[303\].sky_inverter
timestamp 1
transform -1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[304\].sky_inverter
timestamp 1
transform -1 0 17848 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[305\].sky_inverter
timestamp 1
transform 1 0 17848 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[306\].sky_inverter
timestamp 1
transform -1 0 17756 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[307\].sky_inverter
timestamp 1
transform 1 0 17756 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[308\].sky_inverter
timestamp 1
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[309\].sky_inverter
timestamp 1
transform -1 0 17940 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[310\].sky_inverter
timestamp 1
transform 1 0 17940 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[311\].sky_inverter
timestamp 1
transform 1 0 18216 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[312\].sky_inverter
timestamp 1
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[313\].sky_inverter
timestamp 1
transform -1 0 18492 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[314\].sky_inverter
timestamp 1
transform 1 0 18676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[315\].sky_inverter
timestamp 1
transform 1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[316\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[317\].sky_inverter
timestamp 1
transform 1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[318\].sky_inverter
timestamp 1
transform 1 0 19780 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[319\].sky_inverter
timestamp 1
transform 1 0 20056 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[320\].sky_inverter
timestamp 1
transform -1 0 19872 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[321\].sky_inverter
timestamp 1
transform 1 0 19872 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[322\].sky_inverter
timestamp 1
transform 1 0 20148 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[323\].sky_inverter
timestamp 1
transform 1 0 20424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[324\].sky_inverter
timestamp 1
transform 1 0 20700 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[325\].sky_inverter
timestamp 1
transform 1 0 21252 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[326\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[327\].sky_inverter
timestamp 1
transform -1 0 21160 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[328\].sky_inverter
timestamp 1
transform 1 0 21160 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[329\].sky_inverter
timestamp 1
transform 1 0 21436 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[330\].sky_inverter
timestamp 1
transform 1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[331\].sky_inverter
timestamp 1
transform 1 0 21988 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[332\].sky_inverter
timestamp 1
transform 1 0 22264 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[333\].sky_inverter
timestamp 1
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[334\].sky_inverter
timestamp 1
transform 1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[335\].sky_inverter
timestamp 1
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[336\].sky_inverter
timestamp 1
transform 1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[337\].sky_inverter
timestamp 1
transform -1 0 23000 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[338\].sky_inverter
timestamp 1
transform 1 0 22908 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[339\].sky_inverter
timestamp 1
transform 1 0 23828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[340\].sky_inverter
timestamp 1
transform 1 0 24104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[341\].sky_inverter
timestamp 1
transform -1 0 23736 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[342\].sky_inverter
timestamp 1
transform 1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[343\].sky_inverter
timestamp 1
transform 1 0 24656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[344\].sky_inverter
timestamp 1
transform -1 0 24288 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[345\].sky_inverter
timestamp 1
transform 1 0 24288 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[346\].sky_inverter
timestamp 1
transform 1 0 24932 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[347\].sky_inverter
timestamp 1
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[348\].sky_inverter
timestamp 1
transform 1 0 25484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[349\].sky_inverter
timestamp 1
transform -1 0 25300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[350\].sky_inverter
timestamp 1
transform 1 0 25116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[351\].sky_inverter
timestamp 1
transform 1 0 26036 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[352\].sky_inverter
timestamp 1
transform -1 0 26036 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[353\].sky_inverter
timestamp 1
transform 1 0 25944 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[354\].sky_inverter
timestamp 1
transform -1 0 25944 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[355\].sky_inverter
timestamp 1
transform -1 0 25668 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[356\].sky_inverter
timestamp 1
transform 1 0 25852 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[357\].sky_inverter
timestamp 1
transform -1 0 25852 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[358\].sky_inverter
timestamp 1
transform 1 0 26128 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[359\].sky_inverter
timestamp 1
transform 1 0 26404 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[360\].sky_inverter
timestamp 1
transform 1 0 26680 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[361\].sky_inverter
timestamp 1
transform 1 0 26956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[362\].sky_inverter
timestamp 1
transform -1 0 26680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[363\].sky_inverter
timestamp 1
transform 1 0 26680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[364\].sky_inverter
timestamp 1
transform 1 0 26956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[365\].sky_inverter
timestamp 1
transform -1 0 26772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[366\].sky_inverter
timestamp 1
transform 1 0 26772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[367\].sky_inverter
timestamp 1
transform -1 0 26680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[368\].sky_inverter
timestamp 1
transform 1 0 27048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[369\].sky_inverter
timestamp 1
transform -1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[370\].sky_inverter
timestamp 1
transform -1 0 26036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[371\].sky_inverter
timestamp 1
transform -1 0 25760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[372\].sky_inverter
timestamp 1
transform -1 0 25392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[373\].sky_inverter
timestamp 1
transform -1 0 25116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[374\].sky_inverter
timestamp 1
transform 1 0 25300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[375\].sky_inverter
timestamp 1
transform -1 0 25300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[376\].sky_inverter
timestamp 1
transform -1 0 25024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[377\].sky_inverter
timestamp 1
transform -1 0 24748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[378\].sky_inverter
timestamp 1
transform -1 0 24472 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[379\].sky_inverter
timestamp 1
transform 1 0 25024 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[380\].sky_inverter
timestamp 1
transform -1 0 25024 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[381\].sky_inverter
timestamp 1
transform -1 0 24748 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[382\].sky_inverter
timestamp 1
transform -1 0 24472 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[383\].sky_inverter
timestamp 1
transform 1 0 24932 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[384\].sky_inverter
timestamp 1
transform -1 0 24932 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[385\].sky_inverter
timestamp 1
transform -1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[386\].sky_inverter
timestamp 1
transform -1 0 24380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[387\].sky_inverter
timestamp 1
transform -1 0 24104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[388\].sky_inverter
timestamp 1
transform -1 0 23552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[389\].sky_inverter
timestamp 1
transform -1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[390\].sky_inverter
timestamp 1
transform -1 0 23000 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[391\].sky_inverter
timestamp 1
transform -1 0 22724 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[392\].sky_inverter
timestamp 1
transform -1 0 22448 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[393\].sky_inverter
timestamp 1
transform -1 0 22356 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[394\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[395\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[396\].sky_inverter
timestamp 1
transform -1 0 22080 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[397\].sky_inverter
timestamp 1
transform 1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[398\].sky_inverter
timestamp 1
transform 1 0 22080 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[399\].sky_inverter
timestamp 1
transform 1 0 22356 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[400\].sky_inverter
timestamp 1
transform -1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[401\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[402\].sky_inverter
timestamp 1
transform 1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[403\].sky_inverter
timestamp 1
transform 1 0 22080 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[404\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[405\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[406\].sky_inverter
timestamp 1
transform -1 0 22264 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[407\].sky_inverter
timestamp 1
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[408\].sky_inverter
timestamp 1
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[409\].sky_inverter
timestamp 1
transform 1 0 22816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[410\].sky_inverter
timestamp 1
transform 1 0 23092 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[411\].sky_inverter
timestamp 1
transform -1 0 22540 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[412\].sky_inverter
timestamp 1
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[413\].sky_inverter
timestamp 1
transform 1 0 22816 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[414\].sky_inverter
timestamp 1
transform -1 0 22264 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[415\].sky_inverter
timestamp 1
transform 1 0 22080 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[416\].sky_inverter
timestamp 1
transform 1 0 22724 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[417\].sky_inverter
timestamp 1
transform -1 0 22724 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[418\].sky_inverter
timestamp 1
transform -1 0 22448 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[419\].sky_inverter
timestamp 1
transform -1 0 22172 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[420\].sky_inverter
timestamp 1
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[421\].sky_inverter
timestamp 1
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[422\].sky_inverter
timestamp 1
transform -1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[423\].sky_inverter
timestamp 1
transform -1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[424\].sky_inverter
timestamp 1
transform -1 0 20792 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[425\].sky_inverter
timestamp 1
transform -1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[426\].sky_inverter
timestamp 1
transform 1 0 20792 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[427\].sky_inverter
timestamp 1
transform -1 0 20792 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[428\].sky_inverter
timestamp 1
transform -1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[429\].sky_inverter
timestamp 1
transform 1 0 20240 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[430\].sky_inverter
timestamp 1
transform 1 0 20976 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[431\].sky_inverter
timestamp 1
transform -1 0 20976 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[432\].sky_inverter
timestamp 1
transform -1 0 20700 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[433\].sky_inverter
timestamp 1
transform -1 0 20424 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[434\].sky_inverter
timestamp 1
transform -1 0 20148 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[435\].sky_inverter
timestamp 1
transform -1 0 19872 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[436\].sky_inverter
timestamp 1
transform -1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[437\].sky_inverter
timestamp 1
transform -1 0 19320 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[438\].sky_inverter
timestamp 1
transform 1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[439\].sky_inverter
timestamp 1
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[440\].sky_inverter
timestamp 1
transform -1 0 19136 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[441\].sky_inverter
timestamp 1
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[442\].sky_inverter
timestamp 1
transform -1 0 18584 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[443\].sky_inverter
timestamp 1
transform -1 0 18308 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[444\].sky_inverter
timestamp 1
transform -1 0 17480 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[445\].sky_inverter
timestamp 1
transform 1 0 17480 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[446\].sky_inverter
timestamp 1
transform 1 0 17756 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[447\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[448\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[449\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[450\].sky_inverter
timestamp 1
transform -1 0 17664 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[451\].sky_inverter
timestamp 1
transform 1 0 17664 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[452\].sky_inverter
timestamp 1
transform 1 0 17940 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[453\].sky_inverter
timestamp 1
transform 1 0 18216 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[454\].sky_inverter
timestamp 1
transform 1 0 18492 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[455\].sky_inverter
timestamp 1
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[456\].sky_inverter
timestamp 1
transform 1 0 18676 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[457\].sky_inverter
timestamp 1
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[458\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[459\].sky_inverter
timestamp 1
transform 1 0 19504 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[460\].sky_inverter
timestamp 1
transform -1 0 19136 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[461\].sky_inverter
timestamp 1
transform 1 0 19136 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[462\].sky_inverter
timestamp 1
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[463\].sky_inverter
timestamp 1
transform 1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[464\].sky_inverter
timestamp 1
transform -1 0 19320 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[465\].sky_inverter
timestamp 1
transform 1 0 19320 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[466\].sky_inverter
timestamp 1
transform 1 0 19596 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[467\].sky_inverter
timestamp 1
transform -1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[468\].sky_inverter
timestamp 1
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[469\].sky_inverter
timestamp 1
transform 1 0 19228 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[470\].sky_inverter
timestamp 1
transform 1 0 19504 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[471\].sky_inverter
timestamp 1
transform -1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[472\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[473\].sky_inverter
timestamp 1
transform -1 0 19228 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[474\].sky_inverter
timestamp 1
transform -1 0 18952 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[475\].sky_inverter
timestamp 1
transform -1 0 18584 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[476\].sky_inverter
timestamp 1
transform -1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[477\].sky_inverter
timestamp 1
transform -1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[478\].sky_inverter
timestamp 1
transform -1 0 17756 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[479\].sky_inverter
timestamp 1
transform -1 0 17664 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[480\].sky_inverter
timestamp 1
transform 1 0 17664 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[481\].sky_inverter
timestamp 1
transform 1 0 17940 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[482\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[483\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[484\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[485\].sky_inverter
timestamp 1
transform -1 0 17112 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[486\].sky_inverter
timestamp 1
transform -1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[487\].sky_inverter
timestamp 1
transform 1 0 16836 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[488\].sky_inverter
timestamp 1
transform 1 0 17112 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[489\].sky_inverter
timestamp 1
transform 1 0 17388 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[490\].sky_inverter
timestamp 1
transform 1 0 17664 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[491\].sky_inverter
timestamp 1
transform -1 0 17204 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[492\].sky_inverter
timestamp 1
transform 1 0 17204 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[493\].sky_inverter
timestamp 1
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[494\].sky_inverter
timestamp 1
transform 1 0 17756 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[495\].sky_inverter
timestamp 1
transform -1 0 17296 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[496\].sky_inverter
timestamp 1
transform 1 0 17296 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[497\].sky_inverter
timestamp 1
transform 1 0 17572 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[498\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[499\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_250.inv_array\[500\].sky_inverter
timestamp 1
transform 1 0 17480 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[0\].sky_inverter
timestamp 1
transform -1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[1\].sky_inverter
timestamp 1
transform -1 0 14996 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[2\].sky_inverter
timestamp 1
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[3\].sky_inverter
timestamp 1
transform -1 0 14720 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[4\].sky_inverter
timestamp 1
transform 1 0 14720 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[5\].sky_inverter
timestamp 1
transform -1 0 14352 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[6\].sky_inverter
timestamp 1
transform -1 0 14076 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[7\].sky_inverter
timestamp 1
transform 1 0 14352 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[8\].sky_inverter
timestamp 1
transform -1 0 13800 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[9\].sky_inverter
timestamp 1
transform -1 0 13524 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[10\].sky_inverter
timestamp 1
transform -1 0 13248 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[11\].sky_inverter
timestamp 1
transform 1 0 12972 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[12\].sky_inverter
timestamp 1
transform 1 0 13524 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[13\].sky_inverter
timestamp 1
transform -1 0 12972 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[14\].sky_inverter
timestamp 1
transform -1 0 12788 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[15\].sky_inverter
timestamp 1
transform -1 0 12328 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[16\].sky_inverter
timestamp 1
transform 1 0 12328 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[17\].sky_inverter
timestamp 1
transform -1 0 12328 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[18\].sky_inverter
timestamp 1
transform 1 0 12328 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[19\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[20\].sky_inverter
timestamp 1
transform -1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[21\].sky_inverter
timestamp 1
transform -1 0 12880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[22\].sky_inverter
timestamp 1
transform -1 0 12788 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[23\].sky_inverter
timestamp 1
transform 1 0 13524 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[24\].sky_inverter
timestamp 1
transform -1 0 13340 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[25\].sky_inverter
timestamp 1
transform -1 0 13064 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[26\].sky_inverter
timestamp 1
transform 1 0 13524 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[27\].sky_inverter
timestamp 1
transform -1 0 13524 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[28\].sky_inverter
timestamp 1
transform -1 0 12972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[29\].sky_inverter
timestamp 1
transform 1 0 12972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[30\].sky_inverter
timestamp 1
transform -1 0 12696 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[31\].sky_inverter
timestamp 1
transform -1 0 12512 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[32\].sky_inverter
timestamp 1
transform 1 0 12512 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[33\].sky_inverter
timestamp 1
transform -1 0 12236 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[34\].sky_inverter
timestamp 1
transform -1 0 11960 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[35\].sky_inverter
timestamp 1
transform -1 0 11684 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[36\].sky_inverter
timestamp 1
transform -1 0 11408 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[37\].sky_inverter
timestamp 1
transform -1 0 11132 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[38\].sky_inverter
timestamp 1
transform 1 0 11132 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[39\].sky_inverter
timestamp 1
transform -1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[40\].sky_inverter
timestamp 1
transform -1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[41\].sky_inverter
timestamp 1
transform -1 0 10304 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[42\].sky_inverter
timestamp 1
transform -1 0 10028 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[43\].sky_inverter
timestamp 1
transform -1 0 9752 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[44\].sky_inverter
timestamp 1
transform 1 0 9752 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[45\].sky_inverter
timestamp 1
transform -1 0 9476 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[46\].sky_inverter
timestamp 1
transform -1 0 9200 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[47\].sky_inverter
timestamp 1
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[48\].sky_inverter
timestamp 1
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[49\].sky_inverter
timestamp 1
transform -1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[50\].sky_inverter
timestamp 1
transform -1 0 9384 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[51\].sky_inverter
timestamp 1
transform 1 0 9568 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[52\].sky_inverter
timestamp 1
transform -1 0 9292 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[53\].sky_inverter
timestamp 1
transform -1 0 9016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[54\].sky_inverter
timestamp 1
transform 1 0 9016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[55\].sky_inverter
timestamp 1
transform 1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[56\].sky_inverter
timestamp 1
transform -1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[57\].sky_inverter
timestamp 1
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[58\].sky_inverter
timestamp 1
transform -1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[59\].sky_inverter
timestamp 1
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[60\].sky_inverter
timestamp 1
transform -1 0 8924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[61\].sky_inverter
timestamp 1
transform -1 0 8648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[62\].sky_inverter
timestamp 1
transform -1 0 8372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[63\].sky_inverter
timestamp 1
transform -1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[64\].sky_inverter
timestamp 1
transform -1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[65\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[66\].sky_inverter
timestamp 1
transform 1 0 7728 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[67\].sky_inverter
timestamp 1
transform -1 0 7268 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[68\].sky_inverter
timestamp 1
transform -1 0 6900 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[69\].sky_inverter
timestamp 1
transform -1 0 5888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[70\].sky_inverter
timestamp 1
transform -1 0 5612 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[71\].sky_inverter
timestamp 1
transform -1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[72\].sky_inverter
timestamp 1
transform -1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[73\].sky_inverter
timestamp 1
transform -1 0 4784 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[74\].sky_inverter
timestamp 1
transform -1 0 4508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[75\].sky_inverter
timestamp 1
transform -1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[76\].sky_inverter
timestamp 1
transform -1 0 2944 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[77\].sky_inverter
timestamp 1
transform -1 0 2668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[78\].sky_inverter
timestamp 1
transform -1 0 2392 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[79\].sky_inverter
timestamp 1
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[80\].sky_inverter
timestamp 1
transform -1 0 1932 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[81\].sky_inverter
timestamp 1
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[82\].sky_inverter
timestamp 1
transform -1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[83\].sky_inverter
timestamp 1
transform -1 0 2208 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[84\].sky_inverter
timestamp 1
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[85\].sky_inverter
timestamp 1
transform -1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[86\].sky_inverter
timestamp 1
transform -1 0 2208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[87\].sky_inverter
timestamp 1
transform -1 0 2024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[88\].sky_inverter
timestamp 1
transform 1 0 2024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[89\].sky_inverter
timestamp 1
transform 1 0 2852 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[90\].sky_inverter
timestamp 1
transform -1 0 2852 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[91\].sky_inverter
timestamp 1
transform -1 0 2576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[92\].sky_inverter
timestamp 1
transform -1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[93\].sky_inverter
timestamp 1
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[94\].sky_inverter
timestamp 1
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[95\].sky_inverter
timestamp 1
transform -1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[96\].sky_inverter
timestamp 1
transform 1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[97\].sky_inverter
timestamp 1
transform 1 0 3588 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[98\].sky_inverter
timestamp 1
transform -1 0 3588 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[99\].sky_inverter
timestamp 1
transform -1 0 3312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[100\].sky_inverter
timestamp 1
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[101\].sky_inverter
timestamp 1
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[102\].sky_inverter
timestamp 1
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[103\].sky_inverter
timestamp 1
transform 1 0 4048 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[104\].sky_inverter
timestamp 1
transform -1 0 3588 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[105\].sky_inverter
timestamp 1
transform 1 0 3588 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[106\].sky_inverter
timestamp 1
transform 1 0 3864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[107\].sky_inverter
timestamp 1
transform -1 0 3864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[108\].sky_inverter
timestamp 1
transform 1 0 3864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[109\].sky_inverter
timestamp 1
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[110\].sky_inverter
timestamp 1
transform -1 0 3588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[111\].sky_inverter
timestamp 1
transform -1 0 3128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[112\].sky_inverter
timestamp 1
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[113\].sky_inverter
timestamp 1
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[114\].sky_inverter
timestamp 1
transform 1 0 3772 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[115\].sky_inverter
timestamp 1
transform -1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[116\].sky_inverter
timestamp 1
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[117\].sky_inverter
timestamp 1
transform 1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[118\].sky_inverter
timestamp 1
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[119\].sky_inverter
timestamp 1
transform 1 0 4048 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[120\].sky_inverter
timestamp 1
transform -1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[121\].sky_inverter
timestamp 1
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[122\].sky_inverter
timestamp 1
transform 1 0 4692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[123\].sky_inverter
timestamp 1
transform -1 0 4416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[124\].sky_inverter
timestamp 1
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[125\].sky_inverter
timestamp 1
transform 1 0 4508 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[126\].sky_inverter
timestamp 1
transform 1 0 4784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[127\].sky_inverter
timestamp 1
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[128\].sky_inverter
timestamp 1
transform -1 0 5336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[129\].sky_inverter
timestamp 1
transform -1 0 4968 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[130\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[131\].sky_inverter
timestamp 1
transform -1 0 5244 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[132\].sky_inverter
timestamp 1
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[133\].sky_inverter
timestamp 1
transform -1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[134\].sky_inverter
timestamp 1
transform -1 0 5244 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[135\].sky_inverter
timestamp 1
transform 1 0 5244 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[136\].sky_inverter
timestamp 1
transform 1 0 5520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[137\].sky_inverter
timestamp 1
transform -1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[138\].sky_inverter
timestamp 1
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[139\].sky_inverter
timestamp 1
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[140\].sky_inverter
timestamp 1
transform -1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[141\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[142\].sky_inverter
timestamp 1
transform 1 0 6348 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[143\].sky_inverter
timestamp 1
transform 1 0 6624 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[144\].sky_inverter
timestamp 1
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[145\].sky_inverter
timestamp 1
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[146\].sky_inverter
timestamp 1
transform 1 0 7452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[147\].sky_inverter
timestamp 1
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[148\].sky_inverter
timestamp 1
transform -1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[149\].sky_inverter
timestamp 1
transform 1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[150\].sky_inverter
timestamp 1
transform -1 0 8096 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[151\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[152\].sky_inverter
timestamp 1
transform -1 0 7820 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[153\].sky_inverter
timestamp 1
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[154\].sky_inverter
timestamp 1
transform 1 0 8188 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[155\].sky_inverter
timestamp 1
transform -1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[156\].sky_inverter
timestamp 1
transform 1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[157\].sky_inverter
timestamp 1
transform -1 0 8188 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[158\].sky_inverter
timestamp 1
transform -1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[159\].sky_inverter
timestamp 1
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[160\].sky_inverter
timestamp 1
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[161\].sky_inverter
timestamp 1
transform -1 0 8648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[162\].sky_inverter
timestamp 1
transform 1 0 8648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[163\].sky_inverter
timestamp 1
transform 1 0 8924 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[164\].sky_inverter
timestamp 1
transform 1 0 9200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[165\].sky_inverter
timestamp 1
transform 1 0 9476 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[166\].sky_inverter
timestamp 1
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[167\].sky_inverter
timestamp 1
transform 1 0 10028 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[168\].sky_inverter
timestamp 1
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[169\].sky_inverter
timestamp 1
transform 1 0 10580 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[170\].sky_inverter
timestamp 1
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[171\].sky_inverter
timestamp 1
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[172\].sky_inverter
timestamp 1
transform -1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[173\].sky_inverter
timestamp 1
transform 1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[174\].sky_inverter
timestamp 1
transform -1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[175\].sky_inverter
timestamp 1
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[176\].sky_inverter
timestamp 1
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[177\].sky_inverter
timestamp 1
transform 1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[178\].sky_inverter
timestamp 1
transform 1 0 12236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[179\].sky_inverter
timestamp 1
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[180\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[181\].sky_inverter
timestamp 1
transform -1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[182\].sky_inverter
timestamp 1
transform -1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[183\].sky_inverter
timestamp 1
transform 1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[184\].sky_inverter
timestamp 1
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[185\].sky_inverter
timestamp 1
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[186\].sky_inverter
timestamp 1
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[187\].sky_inverter
timestamp 1
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[188\].sky_inverter
timestamp 1
transform 1 0 14444 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[189\].sky_inverter
timestamp 1
transform 1 0 14720 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[190\].sky_inverter
timestamp 1
transform 1 0 15272 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[191\].sky_inverter
timestamp 1
transform -1 0 15272 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[192\].sky_inverter
timestamp 1
transform 1 0 15548 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[193\].sky_inverter
timestamp 1
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[194\].sky_inverter
timestamp 1
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[195\].sky_inverter
timestamp 1
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[196\].sky_inverter
timestamp 1
transform -1 0 15088 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[197\].sky_inverter
timestamp 1
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[198\].sky_inverter
timestamp 1
transform 1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[199\].sky_inverter
timestamp 1
transform 1 0 15640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[200\].sky_inverter
timestamp 1
transform 1 0 15916 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[201\].sky_inverter
timestamp 1
transform -1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[202\].sky_inverter
timestamp 1
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[203\].sky_inverter
timestamp 1
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[204\].sky_inverter
timestamp 1
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[205\].sky_inverter
timestamp 1
transform -1 0 15180 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[206\].sky_inverter
timestamp 1
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[207\].sky_inverter
timestamp 1
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[208\].sky_inverter
timestamp 1
transform 1 0 15732 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[209\].sky_inverter
timestamp 1
transform -1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[210\].sky_inverter
timestamp 1
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[211\].sky_inverter
timestamp 1
transform -1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[212\].sky_inverter
timestamp 1
transform -1 0 14628 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[213\].sky_inverter
timestamp 1
transform -1 0 14352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[214\].sky_inverter
timestamp 1
transform -1 0 14076 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[215\].sky_inverter
timestamp 1
transform -1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[216\].sky_inverter
timestamp 1
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[217\].sky_inverter
timestamp 1
transform -1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[218\].sky_inverter
timestamp 1
transform 1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[219\].sky_inverter
timestamp 1
transform -1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[220\].sky_inverter
timestamp 1
transform -1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[221\].sky_inverter
timestamp 1
transform -1 0 13616 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[222\].sky_inverter
timestamp 1
transform 1 0 13616 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[223\].sky_inverter
timestamp 1
transform -1 0 13340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[224\].sky_inverter
timestamp 1
transform -1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[225\].sky_inverter
timestamp 1
transform -1 0 12788 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[226\].sky_inverter
timestamp 1
transform -1 0 12512 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[227\].sky_inverter
timestamp 1
transform -1 0 12236 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[228\].sky_inverter
timestamp 1
transform -1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[229\].sky_inverter
timestamp 1
transform -1 0 11684 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[230\].sky_inverter
timestamp 1
transform -1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[231\].sky_inverter
timestamp 1
transform 1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[232\].sky_inverter
timestamp 1
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[233\].sky_inverter
timestamp 1
transform -1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[234\].sky_inverter
timestamp 1
transform 1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[235\].sky_inverter
timestamp 1
transform -1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[236\].sky_inverter
timestamp 1
transform -1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[237\].sky_inverter
timestamp 1
transform -1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[238\].sky_inverter
timestamp 1
transform -1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[239\].sky_inverter
timestamp 1
transform -1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[240\].sky_inverter
timestamp 1
transform -1 0 9292 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[241\].sky_inverter
timestamp 1
transform -1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[242\].sky_inverter
timestamp 1
transform 1 0 9016 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[243\].sky_inverter
timestamp 1
transform -1 0 8740 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[244\].sky_inverter
timestamp 1
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[245\].sky_inverter
timestamp 1
transform -1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[246\].sky_inverter
timestamp 1
transform -1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[247\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[248\].sky_inverter
timestamp 1
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[249\].sky_inverter
timestamp 1
transform -1 0 7452 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[250\].sky_inverter
timestamp 1
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[251\].sky_inverter
timestamp 1
transform 1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[252\].sky_inverter
timestamp 1
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[253\].sky_inverter
timestamp 1
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[254\].sky_inverter
timestamp 1
transform -1 0 7452 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[255\].sky_inverter
timestamp 1
transform -1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[256\].sky_inverter
timestamp 1
transform 1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[257\].sky_inverter
timestamp 1
transform -1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[258\].sky_inverter
timestamp 1
transform 1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[259\].sky_inverter
timestamp 1
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[260\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[261\].sky_inverter
timestamp 1
transform 1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[262\].sky_inverter
timestamp 1
transform 1 0 8924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[263\].sky_inverter
timestamp 1
transform 1 0 9200 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[264\].sky_inverter
timestamp 1
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[265\].sky_inverter
timestamp 1
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[266\].sky_inverter
timestamp 1
transform -1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[267\].sky_inverter
timestamp 1
transform 1 0 9936 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[268\].sky_inverter
timestamp 1
transform 1 0 10212 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[269\].sky_inverter
timestamp 1
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[270\].sky_inverter
timestamp 1
transform -1 0 9936 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[271\].sky_inverter
timestamp 1
transform 1 0 10028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[272\].sky_inverter
timestamp 1
transform 1 0 10304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[273\].sky_inverter
timestamp 1
transform -1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[274\].sky_inverter
timestamp 1
transform -1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[275\].sky_inverter
timestamp 1
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[276\].sky_inverter
timestamp 1
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[277\].sky_inverter
timestamp 1
transform 1 0 11500 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[278\].sky_inverter
timestamp 1
transform -1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[279\].sky_inverter
timestamp 1
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[280\].sky_inverter
timestamp 1
transform -1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[281\].sky_inverter
timestamp 1
transform 1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[282\].sky_inverter
timestamp 1
transform 1 0 11776 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[283\].sky_inverter
timestamp 1
transform -1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[284\].sky_inverter
timestamp 1
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[285\].sky_inverter
timestamp 1
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[286\].sky_inverter
timestamp 1
transform 1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[287\].sky_inverter
timestamp 1
transform 1 0 12972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[288\].sky_inverter
timestamp 1
transform -1 0 12972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[289\].sky_inverter
timestamp 1
transform -1 0 12696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[290\].sky_inverter
timestamp 1
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[291\].sky_inverter
timestamp 1
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[292\].sky_inverter
timestamp 1
transform 1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[293\].sky_inverter
timestamp 1
transform 1 0 13524 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[294\].sky_inverter
timestamp 1
transform 1 0 13800 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[295\].sky_inverter
timestamp 1
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[296\].sky_inverter
timestamp 1
transform -1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[297\].sky_inverter
timestamp 1
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[298\].sky_inverter
timestamp 1
transform 1 0 15088 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[299\].sky_inverter
timestamp 1
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[300\].sky_inverter
timestamp 1
transform 1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[301\].sky_inverter
timestamp 1
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[302\].sky_inverter
timestamp 1
transform 1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[303\].sky_inverter
timestamp 1
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[304\].sky_inverter
timestamp 1
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[305\].sky_inverter
timestamp 1
transform 1 0 15640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[306\].sky_inverter
timestamp 1
transform 1 0 15916 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[307\].sky_inverter
timestamp 1
transform 1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[308\].sky_inverter
timestamp 1
transform -1 0 15640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[309\].sky_inverter
timestamp 1
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[310\].sky_inverter
timestamp 1
transform -1 0 15088 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[311\].sky_inverter
timestamp 1
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[312\].sky_inverter
timestamp 1
transform -1 0 14536 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[313\].sky_inverter
timestamp 1
transform -1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[314\].sky_inverter
timestamp 1
transform -1 0 13984 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[315\].sky_inverter
timestamp 1
transform 1 0 13800 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[316\].sky_inverter
timestamp 1
transform -1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[317\].sky_inverter
timestamp 1
transform -1 0 13616 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[318\].sky_inverter
timestamp 1
transform 1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[319\].sky_inverter
timestamp 1
transform -1 0 13156 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[320\].sky_inverter
timestamp 1
transform -1 0 12880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[321\].sky_inverter
timestamp 1
transform -1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[322\].sky_inverter
timestamp 1
transform -1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[323\].sky_inverter
timestamp 1
transform -1 0 12052 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[324\].sky_inverter
timestamp 1
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[325\].sky_inverter
timestamp 1
transform -1 0 11776 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[326\].sky_inverter
timestamp 1
transform -1 0 11500 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[327\].sky_inverter
timestamp 1
transform 1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[328\].sky_inverter
timestamp 1
transform -1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[329\].sky_inverter
timestamp 1
transform -1 0 11132 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[330\].sky_inverter
timestamp 1
transform -1 0 10856 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[331\].sky_inverter
timestamp 1
transform -1 0 10580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[332\].sky_inverter
timestamp 1
transform -1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[333\].sky_inverter
timestamp 1
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[334\].sky_inverter
timestamp 1
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[335\].sky_inverter
timestamp 1
transform -1 0 10120 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[336\].sky_inverter
timestamp 1
transform -1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[337\].sky_inverter
timestamp 1
transform -1 0 9568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[338\].sky_inverter
timestamp 1
transform -1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[339\].sky_inverter
timestamp 1
transform -1 0 9016 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[340\].sky_inverter
timestamp 1
transform -1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[341\].sky_inverter
timestamp 1
transform 1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[342\].sky_inverter
timestamp 1
transform -1 0 8464 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[343\].sky_inverter
timestamp 1
transform -1 0 8280 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[344\].sky_inverter
timestamp 1
transform 1 0 9108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[345\].sky_inverter
timestamp 1
transform -1 0 9108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[346\].sky_inverter
timestamp 1
transform -1 0 8832 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[347\].sky_inverter
timestamp 1
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[348\].sky_inverter
timestamp 1
transform 1 0 9384 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[349\].sky_inverter
timestamp 1
transform -1 0 9384 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[350\].sky_inverter
timestamp 1
transform -1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[351\].sky_inverter
timestamp 1
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[352\].sky_inverter
timestamp 1
transform -1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[353\].sky_inverter
timestamp 1
transform -1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[354\].sky_inverter
timestamp 1
transform 1 0 9476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[355\].sky_inverter
timestamp 1
transform -1 0 9200 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[356\].sky_inverter
timestamp 1
transform -1 0 8924 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[357\].sky_inverter
timestamp 1
transform 1 0 9200 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[358\].sky_inverter
timestamp 1
transform -1 0 8648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[359\].sky_inverter
timestamp 1
transform -1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[360\].sky_inverter
timestamp 1
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[361\].sky_inverter
timestamp 1
transform -1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[362\].sky_inverter
timestamp 1
transform -1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[363\].sky_inverter
timestamp 1
transform -1 0 7636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[364\].sky_inverter
timestamp 1
transform -1 0 7360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[365\].sky_inverter
timestamp 1
transform -1 0 7268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[366\].sky_inverter
timestamp 1
transform -1 0 6992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[367\].sky_inverter
timestamp 1
transform -1 0 6716 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[368\].sky_inverter
timestamp 1
transform -1 0 6532 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[369\].sky_inverter
timestamp 1
transform -1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[370\].sky_inverter
timestamp 1
transform 1 0 6532 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[371\].sky_inverter
timestamp 1
transform -1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[372\].sky_inverter
timestamp 1
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[373\].sky_inverter
timestamp 1
transform -1 0 5704 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[374\].sky_inverter
timestamp 1
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[375\].sky_inverter
timestamp 1
transform -1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[376\].sky_inverter
timestamp 1
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[377\].sky_inverter
timestamp 1
transform 1 0 6992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[378\].sky_inverter
timestamp 1
transform -1 0 6992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[379\].sky_inverter
timestamp 1
transform 1 0 7268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[380\].sky_inverter
timestamp 1
transform -1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[381\].sky_inverter
timestamp 1
transform 1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[382\].sky_inverter
timestamp 1
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[383\].sky_inverter
timestamp 1
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[384\].sky_inverter
timestamp 1
transform -1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[385\].sky_inverter
timestamp 1
transform 1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[386\].sky_inverter
timestamp 1
transform 1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[387\].sky_inverter
timestamp 1
transform -1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[388\].sky_inverter
timestamp 1
transform 1 0 6716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[389\].sky_inverter
timestamp 1
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[390\].sky_inverter
timestamp 1
transform 1 0 7268 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[391\].sky_inverter
timestamp 1
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[392\].sky_inverter
timestamp 1
transform -1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[393\].sky_inverter
timestamp 1
transform -1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[394\].sky_inverter
timestamp 1
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[395\].sky_inverter
timestamp 1
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[396\].sky_inverter
timestamp 1
transform -1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[397\].sky_inverter
timestamp 1
transform 1 0 7544 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[398\].sky_inverter
timestamp 1
transform 1 0 7820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[399\].sky_inverter
timestamp 1
transform 1 0 8096 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[400\].sky_inverter
timestamp 1
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[401\].sky_inverter
timestamp 1
transform 1 0 9292 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[402\].sky_inverter
timestamp 1
transform -1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[403\].sky_inverter
timestamp 1
transform 1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[404\].sky_inverter
timestamp 1
transform -1 0 9108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[405\].sky_inverter
timestamp 1
transform 1 0 9108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[406\].sky_inverter
timestamp 1
transform 1 0 9384 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[407\].sky_inverter
timestamp 1
transform -1 0 8832 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[408\].sky_inverter
timestamp 1
transform 1 0 8648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[409\].sky_inverter
timestamp 1
transform 1 0 8924 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[410\].sky_inverter
timestamp 1
transform 1 0 9476 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[411\].sky_inverter
timestamp 1
transform -1 0 9476 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[412\].sky_inverter
timestamp 1
transform -1 0 9016 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[413\].sky_inverter
timestamp 1
transform 1 0 9016 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[414\].sky_inverter
timestamp 1
transform 1 0 9292 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[415\].sky_inverter
timestamp 1
transform 1 0 9568 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[416\].sky_inverter
timestamp 1
transform 1 0 9844 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[417\].sky_inverter
timestamp 1
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[418\].sky_inverter
timestamp 1
transform -1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[419\].sky_inverter
timestamp 1
transform -1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[420\].sky_inverter
timestamp 1
transform 1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[421\].sky_inverter
timestamp 1
transform 1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[422\].sky_inverter
timestamp 1
transform 1 0 11592 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[423\].sky_inverter
timestamp 1
transform -1 0 11592 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[424\].sky_inverter
timestamp 1
transform -1 0 11316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[425\].sky_inverter
timestamp 1
transform -1 0 10948 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[426\].sky_inverter
timestamp 1
transform 1 0 11776 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[427\].sky_inverter
timestamp 1
transform -1 0 11776 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[428\].sky_inverter
timestamp 1
transform -1 0 11500 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[429\].sky_inverter
timestamp 1
transform -1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[430\].sky_inverter
timestamp 1
transform 1 0 10948 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[431\].sky_inverter
timestamp 1
transform -1 0 10856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[432\].sky_inverter
timestamp 1
transform 1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[433\].sky_inverter
timestamp 1
transform -1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[434\].sky_inverter
timestamp 1
transform -1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[435\].sky_inverter
timestamp 1
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[436\].sky_inverter
timestamp 1
transform 1 0 11684 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[437\].sky_inverter
timestamp 1
transform -1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[438\].sky_inverter
timestamp 1
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[439\].sky_inverter
timestamp 1
transform 1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[440\].sky_inverter
timestamp 1
transform 1 0 12236 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[441\].sky_inverter
timestamp 1
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[442\].sky_inverter
timestamp 1
transform 1 0 12696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[443\].sky_inverter
timestamp 1
transform 1 0 12880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[444\].sky_inverter
timestamp 1
transform 1 0 13248 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[445\].sky_inverter
timestamp 1
transform -1 0 13432 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[446\].sky_inverter
timestamp 1
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[447\].sky_inverter
timestamp 1
transform 1 0 13708 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[448\].sky_inverter
timestamp 1
transform 1 0 13984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[449\].sky_inverter
timestamp 1
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[450\].sky_inverter
timestamp 1
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[451\].sky_inverter
timestamp 1
transform 1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[452\].sky_inverter
timestamp 1
transform -1 0 14352 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[453\].sky_inverter
timestamp 1
transform 1 0 14352 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[454\].sky_inverter
timestamp 1
transform -1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[455\].sky_inverter
timestamp 1
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[456\].sky_inverter
timestamp 1
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[457\].sky_inverter
timestamp 1
transform -1 0 13432 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[458\].sky_inverter
timestamp 1
transform -1 0 13156 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[459\].sky_inverter
timestamp 1
transform -1 0 12880 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[460\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[461\].sky_inverter
timestamp 1
transform 1 0 13432 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[462\].sky_inverter
timestamp 1
transform 1 0 13708 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[463\].sky_inverter
timestamp 1
transform 1 0 13984 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[464\].sky_inverter
timestamp 1
transform -1 0 13432 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[465\].sky_inverter
timestamp 1
transform 1 0 13708 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[466\].sky_inverter
timestamp 1
transform 1 0 13984 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[467\].sky_inverter
timestamp 1
transform 1 0 14260 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[468\].sky_inverter
timestamp 1
transform 1 0 14536 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[469\].sky_inverter
timestamp 1
transform 1 0 14812 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[470\].sky_inverter
timestamp 1
transform 1 0 15088 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[471\].sky_inverter
timestamp 1
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[472\].sky_inverter
timestamp 1
transform -1 0 15732 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[473\].sky_inverter
timestamp 1
transform 1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[474\].sky_inverter
timestamp 1
transform -1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[475\].sky_inverter
timestamp 1
transform -1 0 15824 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[476\].sky_inverter
timestamp 1
transform 1 0 16284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[477\].sky_inverter
timestamp 1
transform -1 0 16284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[478\].sky_inverter
timestamp 1
transform -1 0 16008 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[479\].sky_inverter
timestamp 1
transform -1 0 15732 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[480\].sky_inverter
timestamp 1
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[481\].sky_inverter
timestamp 1
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[482\].sky_inverter
timestamp 1
transform -1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[483\].sky_inverter
timestamp 1
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[484\].sky_inverter
timestamp 1
transform -1 0 15916 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[485\].sky_inverter
timestamp 1
transform 1 0 15916 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[486\].sky_inverter
timestamp 1
transform 1 0 16192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[487\].sky_inverter
timestamp 1
transform 1 0 16468 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[488\].sky_inverter
timestamp 1
transform 1 0 16744 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[489\].sky_inverter
timestamp 1
transform 1 0 17020 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[490\].sky_inverter
timestamp 1
transform 1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[491\].sky_inverter
timestamp 1
transform 1 0 17572 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[492\].sky_inverter
timestamp 1
transform 1 0 18032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[493\].sky_inverter
timestamp 1
transform -1 0 18032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[494\].sky_inverter
timestamp 1
transform -1 0 17756 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[495\].sky_inverter
timestamp 1
transform -1 0 17480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[496\].sky_inverter
timestamp 1
transform 1 0 17940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[497\].sky_inverter
timestamp 1
transform -1 0 17940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[498\].sky_inverter
timestamp 1
transform -1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[499\].sky_inverter
timestamp 1
transform 1 0 17388 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[500\].sky_inverter
timestamp 1
transform 1 0 17664 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[501\].sky_inverter
timestamp 1
transform 1 0 17940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[502\].sky_inverter
timestamp 1
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[503\].sky_inverter
timestamp 1
transform 1 0 18492 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[504\].sky_inverter
timestamp 1
transform 1 0 18768 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[505\].sky_inverter
timestamp 1
transform 1 0 19044 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[506\].sky_inverter
timestamp 1
transform 1 0 19320 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[507\].sky_inverter
timestamp 1
transform 1 0 19596 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[508\].sky_inverter
timestamp 1
transform 1 0 19872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[509\].sky_inverter
timestamp 1
transform -1 0 19688 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[510\].sky_inverter
timestamp 1
transform 1 0 19688 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[511\].sky_inverter
timestamp 1
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[512\].sky_inverter
timestamp 1
transform 1 0 20240 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[513\].sky_inverter
timestamp 1
transform -1 0 20056 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[514\].sky_inverter
timestamp 1
transform 1 0 20056 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[515\].sky_inverter
timestamp 1
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[516\].sky_inverter
timestamp 1
transform -1 0 19780 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[517\].sky_inverter
timestamp 1
transform -1 0 19504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[518\].sky_inverter
timestamp 1
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[519\].sky_inverter
timestamp 1
transform -1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[520\].sky_inverter
timestamp 1
transform -1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[521\].sky_inverter
timestamp 1
transform 1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[522\].sky_inverter
timestamp 1
transform -1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[523\].sky_inverter
timestamp 1
transform 1 0 18768 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[524\].sky_inverter
timestamp 1
transform 1 0 19044 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[525\].sky_inverter
timestamp 1
transform 1 0 19320 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[526\].sky_inverter
timestamp 1
transform -1 0 18768 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[527\].sky_inverter
timestamp 1
transform 1 0 19228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[528\].sky_inverter
timestamp 1
transform -1 0 19228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[529\].sky_inverter
timestamp 1
transform -1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[530\].sky_inverter
timestamp 1
transform -1 0 18492 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[531\].sky_inverter
timestamp 1
transform -1 0 18216 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[532\].sky_inverter
timestamp 1
transform -1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[533\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[534\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[535\].sky_inverter
timestamp 1
transform -1 0 17296 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[536\].sky_inverter
timestamp 1
transform 1 0 17296 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[537\].sky_inverter
timestamp 1
transform 1 0 17572 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[538\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[539\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[540\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[541\].sky_inverter
timestamp 1
transform 1 0 17940 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[542\].sky_inverter
timestamp 1
transform 1 0 18216 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[543\].sky_inverter
timestamp 1
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[544\].sky_inverter
timestamp 1
transform 1 0 18676 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[545\].sky_inverter
timestamp 1
transform 1 0 18952 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[546\].sky_inverter
timestamp 1
transform 1 0 19228 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[547\].sky_inverter
timestamp 1
transform 1 0 19504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[548\].sky_inverter
timestamp 1
transform 1 0 19780 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[549\].sky_inverter
timestamp 1
transform -1 0 19964 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[550\].sky_inverter
timestamp 1
transform 1 0 20056 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[551\].sky_inverter
timestamp 1
transform 1 0 20332 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[552\].sky_inverter
timestamp 1
transform 1 0 20608 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[553\].sky_inverter
timestamp 1
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[554\].sky_inverter
timestamp 1
transform -1 0 20792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[555\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[556\].sky_inverter
timestamp 1
transform -1 0 21528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[557\].sky_inverter
timestamp 1
transform -1 0 21068 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[558\].sky_inverter
timestamp 1
transform 1 0 21344 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[559\].sky_inverter
timestamp 1
transform -1 0 21344 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[560\].sky_inverter
timestamp 1
transform -1 0 21068 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[561\].sky_inverter
timestamp 1
transform -1 0 20792 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[562\].sky_inverter
timestamp 1
transform -1 0 20608 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[563\].sky_inverter
timestamp 1
transform 1 0 21252 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[564\].sky_inverter
timestamp 1
transform -1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[565\].sky_inverter
timestamp 1
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[566\].sky_inverter
timestamp 1
transform 1 0 20700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[567\].sky_inverter
timestamp 1
transform 1 0 20976 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[568\].sky_inverter
timestamp 1
transform 1 0 21252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[569\].sky_inverter
timestamp 1
transform 1 0 21528 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[570\].sky_inverter
timestamp 1
transform 1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[571\].sky_inverter
timestamp 1
transform 1 0 22080 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[572\].sky_inverter
timestamp 1
transform 1 0 22356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[573\].sky_inverter
timestamp 1
transform 1 0 22632 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[574\].sky_inverter
timestamp 1
transform 1 0 22908 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[575\].sky_inverter
timestamp 1
transform 1 0 23184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[576\].sky_inverter
timestamp 1
transform 1 0 23460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[577\].sky_inverter
timestamp 1
transform 1 0 23828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[578\].sky_inverter
timestamp 1
transform 1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[579\].sky_inverter
timestamp 1
transform 1 0 24380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[580\].sky_inverter
timestamp 1
transform -1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[581\].sky_inverter
timestamp 1
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[582\].sky_inverter
timestamp 1
transform 1 0 24288 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[583\].sky_inverter
timestamp 1
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[584\].sky_inverter
timestamp 1
transform 1 0 24840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[585\].sky_inverter
timestamp 1
transform 1 0 25116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[586\].sky_inverter
timestamp 1
transform 1 0 25392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[587\].sky_inverter
timestamp 1
transform 1 0 25668 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[588\].sky_inverter
timestamp 1
transform 1 0 25944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[589\].sky_inverter
timestamp 1
transform 1 0 26404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[590\].sky_inverter
timestamp 1
transform 1 0 26680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[591\].sky_inverter
timestamp 1
transform 1 0 26956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[592\].sky_inverter
timestamp 1
transform -1 0 26588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[593\].sky_inverter
timestamp 1
transform 1 0 27140 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[594\].sky_inverter
timestamp 1
transform -1 0 27140 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[595\].sky_inverter
timestamp 1
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[596\].sky_inverter
timestamp 1
transform 1 0 27508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[597\].sky_inverter
timestamp 1
transform -1 0 27508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[598\].sky_inverter
timestamp 1
transform -1 0 27232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[599\].sky_inverter
timestamp 1
transform -1 0 26956 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[600\].sky_inverter
timestamp 1
transform -1 0 26680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[601\].sky_inverter
timestamp 1
transform 1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[602\].sky_inverter
timestamp 1
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[603\].sky_inverter
timestamp 1
transform -1 0 26588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[604\].sky_inverter
timestamp 1
transform -1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[605\].sky_inverter
timestamp 1
transform -1 0 25392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[606\].sky_inverter
timestamp 1
transform 1 0 25760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[607\].sky_inverter
timestamp 1
transform -1 0 25760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[608\].sky_inverter
timestamp 1
transform -1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[609\].sky_inverter
timestamp 1
transform 1 0 25208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[610\].sky_inverter
timestamp 1
transform -1 0 24564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[611\].sky_inverter
timestamp 1
transform 1 0 24932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[612\].sky_inverter
timestamp 1
transform -1 0 24932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[613\].sky_inverter
timestamp 1
transform -1 0 24656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[614\].sky_inverter
timestamp 1
transform -1 0 24380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[615\].sky_inverter
timestamp 1
transform -1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[616\].sky_inverter
timestamp 1
transform -1 0 23736 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[617\].sky_inverter
timestamp 1
transform -1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[618\].sky_inverter
timestamp 1
transform -1 0 23184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[619\].sky_inverter
timestamp 1
transform -1 0 22908 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[620\].sky_inverter
timestamp 1
transform -1 0 22632 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[621\].sky_inverter
timestamp 1
transform -1 0 22356 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[622\].sky_inverter
timestamp 1
transform -1 0 22080 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[623\].sky_inverter
timestamp 1
transform -1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[624\].sky_inverter
timestamp 1
transform -1 0 21528 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[625\].sky_inverter
timestamp 1
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[626\].sky_inverter
timestamp 1
transform -1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[627\].sky_inverter
timestamp 1
transform -1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[628\].sky_inverter
timestamp 1
transform -1 0 21160 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[629\].sky_inverter
timestamp 1
transform 1 0 21252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[630\].sky_inverter
timestamp 1
transform -1 0 21252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[631\].sky_inverter
timestamp 1
transform -1 0 20976 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[632\].sky_inverter
timestamp 1
transform -1 0 20700 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[633\].sky_inverter
timestamp 1
transform -1 0 20424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[634\].sky_inverter
timestamp 1
transform 1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[635\].sky_inverter
timestamp 1
transform -1 0 20056 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[636\].sky_inverter
timestamp 1
transform 1 0 20424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[637\].sky_inverter
timestamp 1
transform -1 0 20424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[638\].sky_inverter
timestamp 1
transform -1 0 20148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[639\].sky_inverter
timestamp 1
transform -1 0 19872 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[640\].sky_inverter
timestamp 1
transform -1 0 18952 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[641\].sky_inverter
timestamp 1
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[642\].sky_inverter
timestamp 1
transform -1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[643\].sky_inverter
timestamp 1
transform -1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[644\].sky_inverter
timestamp 1
transform -1 0 18768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[645\].sky_inverter
timestamp 1
transform -1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[646\].sky_inverter
timestamp 1
transform -1 0 18216 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[647\].sky_inverter
timestamp 1
transform -1 0 17940 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[648\].sky_inverter
timestamp 1
transform -1 0 17664 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[649\].sky_inverter
timestamp 1
transform -1 0 17388 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[650\].sky_inverter
timestamp 1
transform -1 0 17204 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[651\].sky_inverter
timestamp 1
transform -1 0 16928 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[652\].sky_inverter
timestamp 1
transform -1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[653\].sky_inverter
timestamp 1
transform -1 0 16376 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[654\].sky_inverter
timestamp 1
transform -1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[655\].sky_inverter
timestamp 1
transform 1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[656\].sky_inverter
timestamp 1
transform -1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[657\].sky_inverter
timestamp 1
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[658\].sky_inverter
timestamp 1
transform 1 0 16652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[659\].sky_inverter
timestamp 1
transform -1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[660\].sky_inverter
timestamp 1
transform 1 0 16376 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[661\].sky_inverter
timestamp 1
transform -1 0 16376 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[662\].sky_inverter
timestamp 1
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[663\].sky_inverter
timestamp 1
transform 1 0 16192 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[664\].sky_inverter
timestamp 1
transform 1 0 16468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[665\].sky_inverter
timestamp 1
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[666\].sky_inverter
timestamp 1
transform -1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[667\].sky_inverter
timestamp 1
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[668\].sky_inverter
timestamp 1
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[669\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[670\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[671\].sky_inverter
timestamp 1
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[672\].sky_inverter
timestamp 1
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[673\].sky_inverter
timestamp 1
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[674\].sky_inverter
timestamp 1
transform 1 0 18584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[675\].sky_inverter
timestamp 1
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[676\].sky_inverter
timestamp 1
transform 1 0 19136 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[677\].sky_inverter
timestamp 1
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[678\].sky_inverter
timestamp 1
transform 1 0 19964 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[679\].sky_inverter
timestamp 1
transform -1 0 19964 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[680\].sky_inverter
timestamp 1
transform -1 0 19872 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[681\].sky_inverter
timestamp 1
transform 1 0 20148 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[682\].sky_inverter
timestamp 1
transform -1 0 20148 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[683\].sky_inverter
timestamp 1
transform 1 0 20424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[684\].sky_inverter
timestamp 1
transform -1 0 20424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[685\].sky_inverter
timestamp 1
transform 1 0 20424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[686\].sky_inverter
timestamp 1
transform 1 0 20700 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[687\].sky_inverter
timestamp 1
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[688\].sky_inverter
timestamp 1
transform 1 0 21528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[689\].sky_inverter
timestamp 1
transform 1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[690\].sky_inverter
timestamp 1
transform 1 0 22080 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[691\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[692\].sky_inverter
timestamp 1
transform -1 0 21988 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[693\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[694\].sky_inverter
timestamp 1
transform 1 0 22908 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[695\].sky_inverter
timestamp 1
transform 1 0 23184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[696\].sky_inverter
timestamp 1
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[697\].sky_inverter
timestamp 1
transform 1 0 23460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[698\].sky_inverter
timestamp 1
transform -1 0 23092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[699\].sky_inverter
timestamp 1
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[700\].sky_inverter
timestamp 1
transform 1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[701\].sky_inverter
timestamp 1
transform -1 0 23184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[702\].sky_inverter
timestamp 1
transform 1 0 23184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[703\].sky_inverter
timestamp 1
transform -1 0 22908 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[704\].sky_inverter
timestamp 1
transform -1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[705\].sky_inverter
timestamp 1
transform -1 0 22356 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[706\].sky_inverter
timestamp 1
transform -1 0 22080 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[707\].sky_inverter
timestamp 1
transform -1 0 21988 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[708\].sky_inverter
timestamp 1
transform 1 0 21988 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[709\].sky_inverter
timestamp 1
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[710\].sky_inverter
timestamp 1
transform -1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[711\].sky_inverter
timestamp 1
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[712\].sky_inverter
timestamp 1
transform -1 0 22080 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[713\].sky_inverter
timestamp 1
transform 1 0 22080 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[714\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[715\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[716\].sky_inverter
timestamp 1
transform -1 0 22540 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[717\].sky_inverter
timestamp 1
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[718\].sky_inverter
timestamp 1
transform 1 0 22816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[719\].sky_inverter
timestamp 1
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[720\].sky_inverter
timestamp 1
transform 1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[721\].sky_inverter
timestamp 1
transform 1 0 23828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[722\].sky_inverter
timestamp 1
transform 1 0 24104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[723\].sky_inverter
timestamp 1
transform 1 0 24380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[724\].sky_inverter
timestamp 1
transform 1 0 24656 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[725\].sky_inverter
timestamp 1
transform 1 0 24932 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[726\].sky_inverter
timestamp 1
transform -1 0 24564 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[727\].sky_inverter
timestamp 1
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[728\].sky_inverter
timestamp 1
transform 1 0 25484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[729\].sky_inverter
timestamp 1
transform -1 0 25116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[730\].sky_inverter
timestamp 1
transform 1 0 24932 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[731\].sky_inverter
timestamp 1
transform 1 0 25760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[732\].sky_inverter
timestamp 1
transform -1 0 25760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[733\].sky_inverter
timestamp 1
transform -1 0 25484 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[734\].sky_inverter
timestamp 1
transform 1 0 26036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[735\].sky_inverter
timestamp 1
transform -1 0 26036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[736\].sky_inverter
timestamp 1
transform -1 0 25760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[737\].sky_inverter
timestamp 1
transform -1 0 25484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[738\].sky_inverter
timestamp 1
transform 1 0 26036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[739\].sky_inverter
timestamp 1
transform -1 0 26036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[740\].sky_inverter
timestamp 1
transform -1 0 25760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[741\].sky_inverter
timestamp 1
transform -1 0 25484 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[742\].sky_inverter
timestamp 1
transform 1 0 25760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[743\].sky_inverter
timestamp 1
transform -1 0 25760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[744\].sky_inverter
timestamp 1
transform -1 0 25484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[745\].sky_inverter
timestamp 1
transform 1 0 25944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[746\].sky_inverter
timestamp 1
transform -1 0 25944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[747\].sky_inverter
timestamp 1
transform -1 0 25668 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[748\].sky_inverter
timestamp 1
transform -1 0 25392 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[749\].sky_inverter
timestamp 1
transform -1 0 25116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[750\].sky_inverter
timestamp 1
transform -1 0 24840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[751\].sky_inverter
timestamp 1
transform -1 0 24564 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[752\].sky_inverter
timestamp 1
transform -1 0 24288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[753\].sky_inverter
timestamp 1
transform 1 0 24472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[754\].sky_inverter
timestamp 1
transform -1 0 24472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[755\].sky_inverter
timestamp 1
transform -1 0 24196 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[756\].sky_inverter
timestamp 1
transform 1 0 24472 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[757\].sky_inverter
timestamp 1
transform -1 0 24472 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[758\].sky_inverter
timestamp 1
transform -1 0 24196 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[759\].sky_inverter
timestamp 1
transform -1 0 23920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[760\].sky_inverter
timestamp 1
transform -1 0 23644 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[761\].sky_inverter
timestamp 1
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[762\].sky_inverter
timestamp 1
transform 1 0 23184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[763\].sky_inverter
timestamp 1
transform -1 0 23184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[764\].sky_inverter
timestamp 1
transform -1 0 22908 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[765\].sky_inverter
timestamp 1
transform -1 0 22632 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[766\].sky_inverter
timestamp 1
transform -1 0 22356 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[767\].sky_inverter
timestamp 1
transform 1 0 22632 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[768\].sky_inverter
timestamp 1
transform -1 0 21988 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[769\].sky_inverter
timestamp 1
transform 1 0 22356 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[770\].sky_inverter
timestamp 1
transform -1 0 22356 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[771\].sky_inverter
timestamp 1
transform -1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[772\].sky_inverter
timestamp 1
transform -1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[773\].sky_inverter
timestamp 1
transform -1 0 21528 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[774\].sky_inverter
timestamp 1
transform -1 0 20976 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[775\].sky_inverter
timestamp 1
transform -1 0 20700 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[776\].sky_inverter
timestamp 1
transform -1 0 20424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[777\].sky_inverter
timestamp 1
transform -1 0 20148 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[778\].sky_inverter
timestamp 1
transform -1 0 19872 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[779\].sky_inverter
timestamp 1
transform -1 0 19596 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[780\].sky_inverter
timestamp 1
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[781\].sky_inverter
timestamp 1
transform 1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[782\].sky_inverter
timestamp 1
transform 1 0 19688 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[783\].sky_inverter
timestamp 1
transform -1 0 19136 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[784\].sky_inverter
timestamp 1
transform -1 0 19136 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[785\].sky_inverter
timestamp 1
transform -1 0 19044 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[786\].sky_inverter
timestamp 1
transform -1 0 18768 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[787\].sky_inverter
timestamp 1
transform -1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[788\].sky_inverter
timestamp 1
transform -1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[789\].sky_inverter
timestamp 1
transform -1 0 17940 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[790\].sky_inverter
timestamp 1
transform -1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[791\].sky_inverter
timestamp 1
transform -1 0 17388 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[792\].sky_inverter
timestamp 1
transform -1 0 17112 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[793\].sky_inverter
timestamp 1
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[794\].sky_inverter
timestamp 1
transform -1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[795\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[796\].sky_inverter
timestamp 1
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[797\].sky_inverter
timestamp 1
transform -1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[798\].sky_inverter
timestamp 1
transform -1 0 17572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[799\].sky_inverter
timestamp 1
transform -1 0 17296 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[800\].sky_inverter
timestamp 1
transform 1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[801\].sky_inverter
timestamp 1
transform -1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[802\].sky_inverter
timestamp 1
transform -1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[803\].sky_inverter
timestamp 1
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[804\].sky_inverter
timestamp 1
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[805\].sky_inverter
timestamp 1
transform -1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[806\].sky_inverter
timestamp 1
transform -1 0 16560 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[807\].sky_inverter
timestamp 1
transform 1 0 16744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[808\].sky_inverter
timestamp 1
transform -1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[809\].sky_inverter
timestamp 1
transform -1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[810\].sky_inverter
timestamp 1
transform 1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[811\].sky_inverter
timestamp 1
transform -1 0 15916 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[812\].sky_inverter
timestamp 1
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[813\].sky_inverter
timestamp 1
transform -1 0 15548 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[814\].sky_inverter
timestamp 1
transform -1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[815\].sky_inverter
timestamp 1
transform -1 0 14996 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[816\].sky_inverter
timestamp 1
transform -1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[817\].sky_inverter
timestamp 1
transform -1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[818\].sky_inverter
timestamp 1
transform -1 0 14352 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[819\].sky_inverter
timestamp 1
transform -1 0 13984 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[820\].sky_inverter
timestamp 1
transform -1 0 13432 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[821\].sky_inverter
timestamp 1
transform -1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[822\].sky_inverter
timestamp 1
transform 1 0 13708 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[823\].sky_inverter
timestamp 1
transform -1 0 13708 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[824\].sky_inverter
timestamp 1
transform -1 0 13432 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[825\].sky_inverter
timestamp 1
transform -1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[826\].sky_inverter
timestamp 1
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[827\].sky_inverter
timestamp 1
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[828\].sky_inverter
timestamp 1
transform -1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[829\].sky_inverter
timestamp 1
transform -1 0 13800 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[830\].sky_inverter
timestamp 1
transform -1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[831\].sky_inverter
timestamp 1
transform 1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[832\].sky_inverter
timestamp 1
transform 1 0 13800 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[833\].sky_inverter
timestamp 1
transform -1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[834\].sky_inverter
timestamp 1
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[835\].sky_inverter
timestamp 1
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[836\].sky_inverter
timestamp 1
transform -1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[837\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[838\].sky_inverter
timestamp 1
transform -1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[839\].sky_inverter
timestamp 1
transform -1 0 12512 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[840\].sky_inverter
timestamp 1
transform -1 0 12236 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[841\].sky_inverter
timestamp 1
transform -1 0 11960 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[842\].sky_inverter
timestamp 1
transform 1 0 11776 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[843\].sky_inverter
timestamp 1
transform -1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[844\].sky_inverter
timestamp 1
transform 1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[845\].sky_inverter
timestamp 1
transform -1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[846\].sky_inverter
timestamp 1
transform -1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[847\].sky_inverter
timestamp 1
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[848\].sky_inverter
timestamp 1
transform -1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[849\].sky_inverter
timestamp 1
transform -1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[850\].sky_inverter
timestamp 1
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[851\].sky_inverter
timestamp 1
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[852\].sky_inverter
timestamp 1
transform 1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[853\].sky_inverter
timestamp 1
transform 1 0 12236 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[854\].sky_inverter
timestamp 1
transform -1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[855\].sky_inverter
timestamp 1
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[856\].sky_inverter
timestamp 1
transform 1 0 11776 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[857\].sky_inverter
timestamp 1
transform -1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[858\].sky_inverter
timestamp 1
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[859\].sky_inverter
timestamp 1
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[860\].sky_inverter
timestamp 1
transform -1 0 11592 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[861\].sky_inverter
timestamp 1
transform -1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[862\].sky_inverter
timestamp 1
transform -1 0 11040 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[863\].sky_inverter
timestamp 1
transform -1 0 10764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[864\].sky_inverter
timestamp 1
transform -1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[865\].sky_inverter
timestamp 1
transform -1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[866\].sky_inverter
timestamp 1
transform -1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[867\].sky_inverter
timestamp 1
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[868\].sky_inverter
timestamp 1
transform -1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[869\].sky_inverter
timestamp 1
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[870\].sky_inverter
timestamp 1
transform -1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[871\].sky_inverter
timestamp 1
transform -1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[872\].sky_inverter
timestamp 1
transform -1 0 9568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[873\].sky_inverter
timestamp 1
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[874\].sky_inverter
timestamp 1
transform -1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[875\].sky_inverter
timestamp 1
transform -1 0 10120 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[876\].sky_inverter
timestamp 1
transform -1 0 9844 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[877\].sky_inverter
timestamp 1
transform -1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[878\].sky_inverter
timestamp 1
transform -1 0 9476 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[879\].sky_inverter
timestamp 1
transform 1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[880\].sky_inverter
timestamp 1
transform -1 0 9016 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[881\].sky_inverter
timestamp 1
transform -1 0 8740 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[882\].sky_inverter
timestamp 1
transform -1 0 8464 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[883\].sky_inverter
timestamp 1
transform -1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[884\].sky_inverter
timestamp 1
transform -1 0 7912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[885\].sky_inverter
timestamp 1
transform -1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[886\].sky_inverter
timestamp 1
transform -1 0 7360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[887\].sky_inverter
timestamp 1
transform -1 0 7084 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[888\].sky_inverter
timestamp 1
transform -1 0 6808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[889\].sky_inverter
timestamp 1
transform -1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[890\].sky_inverter
timestamp 1
transform -1 0 6256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[891\].sky_inverter
timestamp 1
transform 1 0 6164 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[892\].sky_inverter
timestamp 1
transform -1 0 6256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[893\].sky_inverter
timestamp 1
transform -1 0 5704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[894\].sky_inverter
timestamp 1
transform -1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[895\].sky_inverter
timestamp 1
transform -1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[896\].sky_inverter
timestamp 1
transform 1 0 4968 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[897\].sky_inverter
timestamp 1
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[898\].sky_inverter
timestamp 1
transform -1 0 4876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[899\].sky_inverter
timestamp 1
transform -1 0 4600 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[900\].sky_inverter
timestamp 1
transform -1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[901\].sky_inverter
timestamp 1
transform 1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[902\].sky_inverter
timestamp 1
transform 1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[903\].sky_inverter
timestamp 1
transform 1 0 4784 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[904\].sky_inverter
timestamp 1
transform -1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[905\].sky_inverter
timestamp 1
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[906\].sky_inverter
timestamp 1
transform 1 0 4232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[907\].sky_inverter
timestamp 1
transform 1 0 4508 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[908\].sky_inverter
timestamp 1
transform 1 0 4784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[909\].sky_inverter
timestamp 1
transform -1 0 4232 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[910\].sky_inverter
timestamp 1
transform 1 0 4232 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[911\].sky_inverter
timestamp 1
transform -1 0 4232 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[912\].sky_inverter
timestamp 1
transform -1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[913\].sky_inverter
timestamp 1
transform 1 0 3956 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[914\].sky_inverter
timestamp 1
transform 1 0 4232 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[915\].sky_inverter
timestamp 1
transform 1 0 4508 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[916\].sky_inverter
timestamp 1
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[917\].sky_inverter
timestamp 1
transform -1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[918\].sky_inverter
timestamp 1
transform -1 0 4324 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[919\].sky_inverter
timestamp 1
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[920\].sky_inverter
timestamp 1
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[921\].sky_inverter
timestamp 1
transform -1 0 4048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[922\].sky_inverter
timestamp 1
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[923\].sky_inverter
timestamp 1
transform 1 0 4508 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[924\].sky_inverter
timestamp 1
transform 1 0 4784 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[925\].sky_inverter
timestamp 1
transform -1 0 4968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[926\].sky_inverter
timestamp 1
transform -1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[927\].sky_inverter
timestamp 1
transform -1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[928\].sky_inverter
timestamp 1
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[929\].sky_inverter
timestamp 1
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[930\].sky_inverter
timestamp 1
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[931\].sky_inverter
timestamp 1
transform -1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[932\].sky_inverter
timestamp 1
transform -1 0 3956 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[933\].sky_inverter
timestamp 1
transform 1 0 3956 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[934\].sky_inverter
timestamp 1
transform 1 0 4232 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[935\].sky_inverter
timestamp 1
transform -1 0 3680 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[936\].sky_inverter
timestamp 1
transform 1 0 3404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[937\].sky_inverter
timestamp 1
transform 1 0 3680 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[938\].sky_inverter
timestamp 1
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[939\].sky_inverter
timestamp 1
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[940\].sky_inverter
timestamp 1
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[941\].sky_inverter
timestamp 1
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[942\].sky_inverter
timestamp 1
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[943\].sky_inverter
timestamp 1
transform 1 0 5060 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[944\].sky_inverter
timestamp 1
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[945\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[946\].sky_inverter
timestamp 1
transform -1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[947\].sky_inverter
timestamp 1
transform 1 0 6532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[948\].sky_inverter
timestamp 1
transform -1 0 6532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[949\].sky_inverter
timestamp 1
transform -1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[950\].sky_inverter
timestamp 1
transform -1 0 5980 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[951\].sky_inverter
timestamp 1
transform -1 0 5704 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[952\].sky_inverter
timestamp 1
transform 1 0 5796 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[953\].sky_inverter
timestamp 1
transform 1 0 6072 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[954\].sky_inverter
timestamp 1
transform 1 0 6348 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[955\].sky_inverter
timestamp 1
transform 1 0 6716 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[956\].sky_inverter
timestamp 1
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[957\].sky_inverter
timestamp 1
transform 1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[958\].sky_inverter
timestamp 1
transform 1 0 7912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[959\].sky_inverter
timestamp 1
transform 1 0 8188 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[960\].sky_inverter
timestamp 1
transform 1 0 8464 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[961\].sky_inverter
timestamp 1
transform 1 0 8740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[962\].sky_inverter
timestamp 1
transform 1 0 9016 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[963\].sky_inverter
timestamp 1
transform 1 0 9568 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[964\].sky_inverter
timestamp 1
transform -1 0 9476 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[965\].sky_inverter
timestamp 1
transform 1 0 9476 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[966\].sky_inverter
timestamp 1
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[967\].sky_inverter
timestamp 1
transform -1 0 10028 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[968\].sky_inverter
timestamp 1
transform 1 0 10028 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[969\].sky_inverter
timestamp 1
transform 1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[970\].sky_inverter
timestamp 1
transform -1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[971\].sky_inverter
timestamp 1
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[972\].sky_inverter
timestamp 1
transform -1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[973\].sky_inverter
timestamp 1
transform -1 0 9384 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[974\].sky_inverter
timestamp 1
transform 1 0 9292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[975\].sky_inverter
timestamp 1
transform -1 0 9292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[976\].sky_inverter
timestamp 1
transform -1 0 9016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[977\].sky_inverter
timestamp 1
transform 1 0 9568 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[978\].sky_inverter
timestamp 1
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[979\].sky_inverter
timestamp 1
transform 1 0 10028 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[980\].sky_inverter
timestamp 1
transform 1 0 10304 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[981\].sky_inverter
timestamp 1
transform 1 0 10488 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[982\].sky_inverter
timestamp 1
transform 1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[983\].sky_inverter
timestamp 1
transform 1 0 11316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[984\].sky_inverter
timestamp 1
transform -1 0 11316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[985\].sky_inverter
timestamp 1
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[986\].sky_inverter
timestamp 1
transform -1 0 11868 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[987\].sky_inverter
timestamp 1
transform -1 0 11316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[988\].sky_inverter
timestamp 1
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[989\].sky_inverter
timestamp 1
transform 1 0 11592 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[990\].sky_inverter
timestamp 1
transform 1 0 12512 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[991\].sky_inverter
timestamp 1
transform -1 0 12236 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[992\].sky_inverter
timestamp 1
transform 1 0 12236 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[993\].sky_inverter
timestamp 1
transform 1 0 12328 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[994\].sky_inverter
timestamp 1
transform 1 0 12604 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[995\].sky_inverter
timestamp 1
transform 1 0 12880 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[996\].sky_inverter
timestamp 1
transform 1 0 13156 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[997\].sky_inverter
timestamp 1
transform 1 0 13524 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[998\].sky_inverter
timestamp 1
transform 1 0 13892 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[999\].sky_inverter
timestamp 1
transform 1 0 14260 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ring_1001.inv_array\[1000\].sky_inverter
timestamp 1
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_19
timestamp 1
transform -1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_20
timestamp 1
transform -1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_21
timestamp 1
transform -1 0 9200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_22
timestamp 1
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_23
timestamp 1
transform -1 0 8096 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_24
timestamp 1
transform -1 0 7544 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_25
timestamp 1
transform -1 0 6992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_26
timestamp 1
transform -1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_27
timestamp 1
transform -1 0 14720 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_28
timestamp 1
transform -1 0 14168 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_29
timestamp 1
transform -1 0 13800 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_30
timestamp 1
transform -1 0 13064 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_31
timestamp 1
transform -1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_32
timestamp 1
transform -1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_33
timestamp 1
transform -1 0 11408 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_34
timestamp 1
transform -1 0 10856 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_35
timestamp 1
transform -1 0 17204 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_36
timestamp 1
transform -1 0 16376 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_tt09_ring_osc_37
timestamp 1
transform -1 0 15916 0 1 21216
box -38 -48 314 592
<< labels >>
flabel metal4 s 4316 496 4636 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12090 496 12410 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19864 496 20184 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27638 496 27958 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11430 496 11750 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19204 496 19524 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26978 496 27298 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
